  --------------------------------------------------------------------------------------------------------------------------
-- Original Authors : Simon Doherty, Eric Lunty, Kyle Brooks, Peter Roland						--
-- Date created: N/A 													--
--															--
-- Additional Authors : Randi Derbyshire, Adam Narten, Oliver Rarog, Celeste Chiasson					--
-- Date edited: March 26, 2018											--
--															--
-- This program takes a value from the synthesizer.vhd file and runs it through the 12-bit ROM to find the 	 	--
-- respective sine wave value. 												--
--------------------------------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use IEEE.STD_LOGIC_SIGNED.all;
use ieee.numeric_std.all;               -- Needed for shifts

entity ClarinetSin_lut is

port (
	clk      : in  std_logic;
	en       : in  std_logic;
	
	--Address input
	address_reg : in std_logic_vector(11 downto 0); 
	
	--Sine value output
	sin_out  : out std_logic_vector(31 downto 0)
	);
end entity;


architecture rtl of ClarinetSin_lut is


type rom_type is array (0 to 4095) of std_logic_vector (11 downto 0);

constant SIN_ROM : rom_type :=

(
X"000", X"02F", X"05E", X"089", X"0B9", X"0E8", X"117", X"142", 
X"171", X"1A0", X"1CF", X"1FA", X"229", X"257", X"286", X"2B0", 
X"2DF", X"30D", X"33B", X"369", X"393", X"3C1", X"3EE", X"41C", 
X"445", X"472", X"49F", X"4CB", X"4F4", X"520", X"54C", X"578", 
X"5A3", X"5CB", X"5F6", X"621", X"64B", X"672", X"69C", X"6C6", 
X"6EF", X"715", X"73E", X"766", X"78F", X"7B3", X"7DB", X"802", 
X"829", X"850", X"872", X"898", X"8BE", X"8E3", X"905", X"929", 
X"94E", X"971", X"992", X"9B5", X"9D7", X"9F9", X"A1B", X"A3A", 
X"A5B", X"A7B", X"A9B", X"AB8", X"AD8", X"AF7", X"B15", X"B30", 
X"B4E", X"B6B", X"B88", X"BA2", X"BBE", X"BD9", X"BF4", X"C0E", 
X"C26", X"C3F", X"C59", X"C71", X"C87", X"C9F", X"CB6", X"CCD", 
X"CE1", X"CF7", X"D0C", X"D21", X"D35", X"D47", X"D5B", X"D6E", 
X"D80", X"D90", X"DA2", X"DB3", X"DC3", X"DD2", X"DE1", X"DF0", 
X"DFF", X"E0C", X"E19", X"E26", X"E33", X"E3F", X"E4A", X"E55", 
X"E5F", X"E6A", X"E73", X"E7C", X"E85", X"E8D", X"E94", X"E9C", 
X"EA3", X"EA9", X"EAF", X"EB4", X"EB9", X"EBE", X"EC2", X"EC6", 
X"EC9", X"ECC", X"ECF", X"ED1", X"ED2", X"ED3", X"ED4", X"ED5", 
X"ED5", X"ED4", X"ED3", X"ED2", X"ED1", X"ECE", X"ECC", X"EC9", 
X"EC6", X"EC3", X"EBF", X"EBA", X"EB6", X"EB1", X"EAC", X"EA6", 
X"EA0", X"E9A", X"E93", X"E8C", X"E85", X"E7E", X"E76", X"E6D", 
X"E65", X"E5D", X"E53", X"E4A", X"E40", X"E37", X"E2D", X"E22", 
X"E17", X"E0C", X"E01", X"DF6", X"DEA", X"DDE", X"DD3", X"DC6", 
X"DB9", X"DAC", X"DA0", X"D93", X"D85", X"D78", X"D6A", X"D5D", 
X"D4F", X"D40", X"D32", X"D24", X"D15", X"D06", X"CF7", X"CE9", 
X"CDA", X"CCA", X"CBB", X"CAC", X"C9C", X"C8C", X"C7C", X"C6C", 
X"C5E", X"C4D", X"C3D", X"C2D", X"C1E", X"C0D", X"BFD", X"BEC", 
X"BDD", X"BCD", X"BBC", X"BAB", X"B9B", X"B8C", X"B7B", X"B6A", 
X"B5A", X"B4B", X"B3A", X"B29", X"B19", X"B0A", X"AF9", X"AE9", 
X"AD9", X"ACA", X"ABA", X"AAA", X"A99", X"A89", X"A7B", X"A6B", 
X"A5B", X"A4C", X"A3D", X"A2E", X"A1F", X"A0F", X"A02", X"9F3", 
X"9E4", X"9D5", X"9C6", X"9B9", X"9AA", X"99C", X"98E", X"981", 
X"973", X"966", X"958", X"94C", X"93F", X"932", X"925", X"919", 
X"90D", X"900", X"8F4", X"8E8", X"8DD", X"8D1", X"8C6", X"8BB", 
X"8B0", X"8A6", X"89B", X"890", X"887", X"87C", X"872", X"869", 
X"85F", X"857", X"84D", X"844", X"83B", X"834", X"82B", X"823", 
X"81B", X"814", X"80C", X"805", X"7FE", X"7F7", X"7F1", X"7EA", 
X"7E4", X"7DE", X"7D8", X"7D2", X"7CD", X"7C8", X"7C3", X"7BE", 
X"7B9", X"7B5", X"7B1", X"7AD", X"7A9", X"7A5", X"7A2", X"79E", 
X"79B", X"798", X"796", X"793", X"791", X"78F", X"78D", X"78B", 
X"78A", X"788", X"787", X"786", X"785", X"784", X"784", X"783", 
X"783", X"783", X"783", X"784", X"784", X"785", X"785", X"786", 
X"787", X"789", X"78A", X"78B", X"78D", X"78F", X"791", X"793", 
X"795", X"797", X"799", X"79C", X"79F", X"7A1", X"7A4", X"7A7", 
X"7AA", X"7AD", X"7B1", X"7B4", X"7B8", X"7BC", X"7BF", X"7C3", 
X"7C7", X"7CB", X"7CE", X"7D3", X"7D7", X"7DB", X"7DF", X"7E4", 
X"7E8", X"7ED", X"7F2", X"7F6", X"7FB", X"7FF", X"804", X"809", 
X"80E", X"813", X"818", X"81C", X"821", X"826", X"82B", X"830", 
X"835", X"83A", X"840", X"845", X"84A", X"84F", X"854", X"859", 
X"85E", X"863", X"868", X"86E", X"872", X"877", X"87C", X"882", 
X"887", X"88B", X"890", X"895", X"89A", X"89F", X"8A4", X"8A9", 
X"8AD", X"8B2", X"8B6", X"8BB", X"8C0", X"8C4", X"8C8", X"8CD", 
X"8D1", X"8D6", X"8DA", X"8DE", X"8E2", X"8E6", X"8EA", X"8EE", 
X"8F2", X"8F5", X"8F9", X"8FC", X"900", X"904", X"907", X"90A", 
X"90D", X"911", X"914", X"916", X"919", X"91C", X"91F", X"922", 
X"924", X"927", X"929", X"92B", X"92D", X"930", X"932", X"934", 
X"935", X"937", X"939", X"93A", X"93C", X"93D", X"93E", X"940", 
X"941", X"942", X"942", X"943", X"944", X"945", X"945", X"945", 
X"946", X"946", X"946", X"946", X"946", X"946", X"946", X"945", 
X"945", X"944", X"944", X"943", X"942", X"941", X"941", X"93F", 
X"93E", X"93D", X"93C", X"93A", X"939", X"937", X"936", X"934", 
X"932", X"930", X"92E", X"92C", X"92A", X"928", X"925", X"923", 
X"921", X"91E", X"91B", X"919", X"916", X"913", X"910", X"90D", 
X"90A", X"907", X"904", X"901", X"8FE", X"8FA", X"8F7", X"8F3", 
X"8F0", X"8EC", X"8E9", X"8E5", X"8E1", X"8DD", X"8D9", X"8D5", 
X"8D1", X"8CE", X"8C9", X"8C5", X"8C1", X"8BD", X"8B9", X"8B4", 
X"8B0", X"8AC", X"8A7", X"8A3", X"89E", X"89A", X"895", X"891", 
X"88C", X"887", X"883", X"87E", X"879", X"874", X"86F", X"86B", 
X"866", X"860", X"85C", X"857", X"852", X"84D", X"848", X"843", 
X"83E", X"838", X"833", X"82E", X"829", X"824", X"81E", X"81A", 
X"814", X"80F", X"809", X"805", X"7FF", X"7FA", X"7F4", X"7EF", 
X"7EA", X"7E4", X"7DF", X"7D9", X"7D4", X"7CF", X"7C9", X"7C4", 
X"7BF", X"7B9", X"7B3", X"7AE", X"7A9", X"7A3", X"79D", X"798", 
X"792", X"78D", X"787", X"782", X"77C", X"777", X"771", X"76B", 
X"766", X"760", X"75B", X"755", X"74F", X"749", X"744", X"73E", 
X"738", X"733", X"72D", X"727", X"722", X"71C", X"716", X"710", 
X"70A", X"704", X"6FF", X"6F9", X"6F3", X"6ED", X"6E7", X"6E1", 
X"6DB", X"6D5", X"6CF", X"6CA", X"6C3", X"6BD", X"6B7", X"6B1", 
X"6AB", X"6A5", X"69F", X"698", X"693", X"68C", X"686", X"67F", 
X"679", X"673", X"66C", X"666", X"660", X"659", X"653", X"64C", 
X"646", X"63F", X"638", X"632", X"62B", X"625", X"61E", X"617", 
X"610", X"609", X"602", X"5FB", X"5F4", X"5EE", X"5E6", X"5DF", 
X"5D8", X"5D1", X"5CA", X"5C2", X"5BB", X"5B3", X"5AD", X"5A5", 
X"59D", X"596", X"58F", X"587", X"57F", X"577", X"570", X"568", 
X"560", X"558", X"550", X"549", X"541", X"539", X"530", X"529", 
X"520", X"518", X"510", X"508", X"4FF", X"4F7", X"4EE", X"4E6", 
X"4DE", X"4D5", X"4CC", X"4C3", X"4BB", X"4B3", X"4AA", X"4A1", 
X"499", X"48F", X"486", X"47D", X"475", X"46C", X"463", X"459", 
X"450", X"448", X"43E", X"435", X"42B", X"423", X"419", X"410", 
X"406", X"3FE", X"3F4", X"3EB", X"3E1", X"3D7", X"3CF", X"3C5", 
X"3BB", X"3B2", X"3A9", X"39F", X"396", X"38C", X"383", X"379", 
X"370", X"366", X"35D", X"353", X"34A", X"340", X"336", X"32D", 
X"324", X"31A", X"310", X"308", X"2FE", X"2F4", X"2EB", X"2E2", 
X"2D9", X"2CF", X"2C6", X"2BC", X"2B4", X"2AB", X"2A1", X"298", 
X"290", X"286", X"27D", X"274", X"26C", X"263", X"25A", X"251", 
X"249", X"241", X"238", X"22F", X"227", X"21F", X"217", X"20F", 
X"207", X"1FF", X"1F7", X"1EF", X"1E7", X"1E0", X"1D9", X"1D1", 
X"1CA", X"1C2", X"1BC", X"1B5", X"1AE", X"1A7", X"1A1", X"19A", 
X"193", X"18D", X"187", X"181", X"17B", X"175", X"170", X"16A", 
X"165", X"15F", X"15A", X"155", X"150", X"14C", X"147", X"143", 
X"13E", X"13A", X"136", X"133", X"12F", X"12C", X"128", X"125", 
X"122", X"11F", X"11D", X"11A", X"118", X"116", X"114", X"112", 
X"111", X"10F", X"10E", X"10D", X"10C", X"10C", X"10B", X"10B", 
X"10B", X"10B", X"10B", X"10C", X"10D", X"10D", X"10F", X"110", 
X"111", X"113", X"115", X"117", X"119", X"11C", X"11F", X"122", 
X"125", X"128", X"12B", X"12F", X"133", X"137", X"13B", X"140", 
X"145", X"14A", X"14F", X"154", X"15A", X"160", X"166", X"16C", 
X"172", X"179", X"180", X"186", X"18E", X"195", X"19D", X"1A4", 
X"1AC", X"1B5", X"1BD", X"1C6", X"1CE", X"1D7", X"1E1", X"1EA", 
X"1F3", X"1FD", X"207", X"211", X"21B", X"225", X"230", X"23B", 
X"245", X"251", X"25C", X"268", X"274", X"27F", X"28B", X"297", 
X"2A4", X"2AF", X"2BC", X"2C9", X"2D6", X"2E2", X"2F0", X"2FD", 
X"30B", X"319", X"326", X"334", X"342", X"350", X"35E", X"36C", 
X"37B", X"38A", X"397", X"3A6", X"3B6", X"3C5", X"3D3", X"3E2", 
X"3F2", X"401", X"411", X"41F", X"42F", X"43F", X"44F", X"45E", 
X"46E", X"47E", X"48E", X"49D", X"4AD", X"4BE", X"4CE", X"4DE", 
X"4ED", X"4FE", X"50E", X"51F", X"52E", X"53E", X"54F", X"55F", 
X"56E", X"57F", X"58F", X"5A0", X"5AF", X"5BF", X"5D0", X"5E0", 
X"5F1", X"5FF", X"610", X"620", X"630", X"63F", X"64F", X"65F", 
X"66F", X"67D", X"68D", X"69C", X"6AC", X"6BC", X"6CA", X"6D9", 
X"6E8", X"6F7", X"705", X"714", X"723", X"731", X"73F", X"74D", 
X"75B", X"769", X"776", X"784", X"792", X"79F", X"7AD", X"7B9", 
X"7C6", X"7D3", X"7E0", X"7EB", X"7F7", X"804", X"810", X"81B", 
X"826", X"832", X"83D", X"848", X"852", X"85D", X"867", X"872", 
X"87B", X"885", X"88E", X"898", X"8A0", X"8A9", X"8B2", X"8BB", 
X"8C2", X"8CA", X"8D2", X"8DA", X"8E1", X"8E8", X"8EE", X"8F5", 
X"8FB", X"901", X"907", X"90D", X"912", X"917", X"91C", X"920", 
X"925", X"929", X"92C", X"930", X"933", X"936", X"939", X"93B", 
X"93E", X"940", X"941", X"943", X"944", X"945", X"945", X"946", 
X"946", X"946", X"945", X"945", X"944", X"943", X"941", X"940", 
X"93E", X"93B", X"939", X"936", X"933", X"930", X"92C", X"929", 
X"925", X"920", X"91C", X"917", X"912", X"90D", X"907", X"901", 
X"8FB", X"8F5", X"8EE", X"8E8", X"8E1", X"8DA", X"8D2", X"8CA", 
X"8C2", X"8BB", X"8B2", X"8A9", X"8A0", X"898", X"88E", X"885", 
X"87B", X"872", X"867", X"85D", X"852", X"848", X"83D", X"832", 
X"826", X"81B", X"810", X"804", X"7F7", X"7EB", X"7E0", X"7D3", 
X"7C6", X"7B9", X"7AD", X"79F", X"792", X"784", X"776", X"769", 
X"75B", X"74D", X"73F", X"731", X"723", X"714", X"705", X"6F7", 
X"6E8", X"6D9", X"6CA", X"6BC", X"6AC", X"69C", X"68D", X"67D", 
X"66F", X"65F", X"64F", X"63F", X"630", X"620", X"610", X"5FF", 
X"5F1", X"5E0", X"5D0", X"5BF", X"5AF", X"5A0", X"58F", X"57F", 
X"56E", X"55F", X"54F", X"53E", X"52E", X"51F", X"50E", X"4FE", 
X"4ED", X"4DE", X"4CE", X"4BE", X"4AD", X"49D", X"48E", X"47E", 
X"46E", X"45E", X"44F", X"43F", X"42F", X"41F", X"411", X"401", 
X"3F2", X"3E2", X"3D3", X"3C5", X"3B6", X"3A6", X"397", X"38A", 
X"37B", X"36C", X"35E", X"350", X"342", X"334", X"326", X"319", 
X"30B", X"2FD", X"2F0", X"2E2", X"2D6", X"2C9", X"2BC", X"2AF", 
X"2A4", X"297", X"28B", X"27F", X"274", X"268", X"25C", X"251", 
X"245", X"23B", X"230", X"225", X"21B", X"211", X"207", X"1FD", 
X"1F3", X"1EA", X"1E1", X"1D7", X"1CE", X"1C6", X"1BD", X"1B5", 
X"1AC", X"1A4", X"19D", X"195", X"18E", X"186", X"180", X"179", 
X"172", X"16C", X"166", X"160", X"15A", X"154", X"14F", X"14A", 
X"145", X"140", X"13B", X"137", X"133", X"12F", X"12B", X"128", 
X"125", X"122", X"11F", X"11C", X"119", X"117", X"115", X"113", 
X"111", X"110", X"10F", X"10D", X"10D", X"10C", X"10B", X"10B", 
X"10B", X"10B", X"10B", X"10C", X"10C", X"10D", X"10E", X"10F", 
X"111", X"112", X"114", X"116", X"118", X"11A", X"11D", X"11F", 
X"122", X"125", X"128", X"12C", X"12F", X"133", X"136", X"13A", 
X"13E", X"143", X"147", X"14C", X"150", X"155", X"15A", X"15F", 
X"165", X"16A", X"170", X"175", X"17B", X"181", X"187", X"18D", 
X"193", X"19A", X"1A1", X"1A7", X"1AE", X"1B5", X"1BC", X"1C2", 
X"1CA", X"1D1", X"1D9", X"1E0", X"1E7", X"1EF", X"1F7", X"1FF", 
X"207", X"20F", X"217", X"21F", X"227", X"22F", X"238", X"241", 
X"249", X"251", X"25A", X"263", X"26C", X"274", X"27D", X"286", 
X"290", X"298", X"2A1", X"2AB", X"2B4", X"2BC", X"2C6", X"2CF", 
X"2D9", X"2E2", X"2EB", X"2F4", X"2FE", X"308", X"310", X"31A", 
X"324", X"32D", X"336", X"340", X"34A", X"353", X"35D", X"366", 
X"370", X"379", X"383", X"38C", X"396", X"39F", X"3A9", X"3B2", 
X"3BB", X"3C5", X"3CF", X"3D7", X"3E1", X"3EB", X"3F4", X"3FE", 
X"406", X"410", X"419", X"423", X"42B", X"435", X"43E", X"448", 
X"450", X"459", X"463", X"46C", X"475", X"47D", X"486", X"48F", 
X"499", X"4A1", X"4AA", X"4B3", X"4BB", X"4C3", X"4CC", X"4D5", 
X"4DE", X"4E6", X"4EE", X"4F7", X"4FF", X"508", X"510", X"518", 
X"520", X"529", X"530", X"539", X"541", X"549", X"550", X"558", 
X"560", X"568", X"570", X"577", X"57F", X"587", X"58F", X"596", 
X"59D", X"5A5", X"5AD", X"5B3", X"5BB", X"5C2", X"5CA", X"5D1", 
X"5D8", X"5DF", X"5E6", X"5EE", X"5F4", X"5FB", X"602", X"609", 
X"610", X"617", X"61E", X"625", X"62B", X"632", X"638", X"63F", 
X"646", X"64C", X"653", X"659", X"660", X"666", X"66C", X"673", 
X"679", X"67F", X"686", X"68C", X"693", X"698", X"69F", X"6A5", 
X"6AB", X"6B1", X"6B7", X"6BD", X"6C3", X"6CA", X"6CF", X"6D5", 
X"6DB", X"6E1", X"6E7", X"6ED", X"6F3", X"6F9", X"6FF", X"704", 
X"70A", X"710", X"716", X"71C", X"722", X"727", X"72D", X"733", 
X"738", X"73E", X"744", X"749", X"74F", X"755", X"75B", X"760", 
X"766", X"76B", X"771", X"777", X"77C", X"782", X"787", X"78D", 
X"792", X"798", X"79D", X"7A3", X"7A9", X"7AE", X"7B3", X"7B9", 
X"7BF", X"7C4", X"7C9", X"7CF", X"7D4", X"7D9", X"7DF", X"7E4", 
X"7EA", X"7EF", X"7F4", X"7FA", X"7FF", X"805", X"809", X"80F", 
X"814", X"81A", X"81E", X"824", X"829", X"82E", X"833", X"838", 
X"83E", X"843", X"848", X"84D", X"852", X"857", X"85C", X"860", 
X"866", X"86B", X"86F", X"874", X"879", X"87E", X"883", X"887", 
X"88C", X"891", X"895", X"89A", X"89E", X"8A3", X"8A7", X"8AC", 
X"8B0", X"8B4", X"8B9", X"8BD", X"8C1", X"8C5", X"8C9", X"8CE", 
X"8D2", X"8D5", X"8D9", X"8DD", X"8E1", X"8E5", X"8E9", X"8EC", 
X"8F0", X"8F3", X"8F7", X"8FA", X"8FE", X"901", X"904", X"907", 
X"90A", X"90D", X"910", X"913", X"916", X"919", X"91B", X"91E", 
X"921", X"923", X"925", X"928", X"92A", X"92C", X"92E", X"930", 
X"932", X"934", X"936", X"937", X"939", X"93A", X"93C", X"93D", 
X"93E", X"93F", X"941", X"941", X"942", X"943", X"944", X"944", 
X"945", X"945", X"946", X"946", X"946", X"946", X"946", X"946", 
X"946", X"945", X"945", X"945", X"944", X"943", X"942", X"942", 
X"941", X"940", X"93E", X"93D", X"93C", X"93A", X"939", X"937", 
X"935", X"934", X"932", X"930", X"92D", X"92B", X"929", X"927", 
X"924", X"922", X"91F", X"91C", X"919", X"916", X"914", X"911", 
X"90D", X"90A", X"907", X"904", X"900", X"8FC", X"8F9", X"8F5", 
X"8F2", X"8EE", X"8EA", X"8E6", X"8E2", X"8DE", X"8DA", X"8D6", 
X"8D1", X"8CD", X"8C8", X"8C4", X"8C0", X"8BB", X"8B6", X"8B2", 
X"8AD", X"8A9", X"8A4", X"89F", X"89A", X"895", X"890", X"88B", 
X"887", X"882", X"87C", X"877", X"872", X"86E", X"868", X"863", 
X"85E", X"859", X"854", X"84F", X"84A", X"845", X"840", X"83A", 
X"835", X"830", X"82B", X"826", X"821", X"81C", X"818", X"813", 
X"80E", X"809", X"804", X"7FF", X"7FB", X"7F6", X"7F2", X"7ED", 
X"7E8", X"7E4", X"7DF", X"7DB", X"7D7", X"7D3", X"7CE", X"7CB", 
X"7C7", X"7C3", X"7BF", X"7BC", X"7B8", X"7B4", X"7B1", X"7AD", 
X"7AA", X"7A7", X"7A4", X"7A1", X"79F", X"79C", X"799", X"797", 
X"795", X"793", X"791", X"78F", X"78D", X"78B", X"78A", X"789", 
X"787", X"786", X"785", X"785", X"784", X"784", X"783", X"783", 
X"783", X"783", X"784", X"784", X"785", X"786", X"787", X"788", 
X"78A", X"78B", X"78D", X"78F", X"791", X"793", X"796", X"798", 
X"79B", X"79E", X"7A2", X"7A5", X"7A9", X"7AD", X"7B1", X"7B5", 
X"7B9", X"7BE", X"7C3", X"7C8", X"7CD", X"7D2", X"7D8", X"7DE", 
X"7E4", X"7EA", X"7F1", X"7F7", X"7FE", X"805", X"80C", X"814", 
X"81B", X"823", X"82B", X"834", X"83B", X"844", X"84D", X"857", 
X"85F", X"869", X"872", X"87C", X"887", X"890", X"89B", X"8A6", 
X"8B0", X"8BB", X"8C6", X"8D1", X"8DD", X"8E8", X"8F4", X"900", 
X"90D", X"919", X"925", X"932", X"93F", X"94C", X"958", X"966", 
X"973", X"981", X"98E", X"99C", X"9AA", X"9B9", X"9C6", X"9D5", 
X"9E4", X"9F3", X"A02", X"A0F", X"A1F", X"A2E", X"A3D", X"A4C", 
X"A5B", X"A6B", X"A7B", X"A89", X"A99", X"AAA", X"ABA", X"ACA", 
X"AD9", X"AE9", X"AF9", X"B0A", X"B19", X"B29", X"B3A", X"B4B", 
X"B5A", X"B6A", X"B7B", X"B8C", X"B9B", X"BAB", X"BBC", X"BCD", 
X"BDD", X"BEC", X"BFD", X"C0D", X"C1E", X"C2D", X"C3D", X"C4D", 
X"C5E", X"C6C", X"C7C", X"C8C", X"C9C", X"CAC", X"CBB", X"CCA", 
X"CDA", X"CE9", X"CF7", X"D06", X"D15", X"D24", X"D32", X"D40", 
X"D4F", X"D5D", X"D6A", X"D78", X"D85", X"D93", X"DA0", X"DAC", 
X"DB9", X"DC6", X"DD3", X"DDE", X"DEA", X"DF6", X"E01", X"E0C", 
X"E17", X"E22", X"E2D", X"E37", X"E40", X"E4A", X"E53", X"E5D", 
X"E65", X"E6D", X"E76", X"E7E", X"E85", X"E8C", X"E93", X"E9A", 
X"EA0", X"EA6", X"EAC", X"EB1", X"EB6", X"EBA", X"EBF", X"EC3", 
X"EC6", X"EC9", X"ECC", X"ECE", X"ED1", X"ED2", X"ED3", X"ED4", 
X"ED5", X"ED5", X"ED4", X"ED3", X"ED2", X"ED1", X"ECF", X"ECC", 
X"EC9", X"EC6", X"EC2", X"EBE", X"EB9", X"EB4", X"EAF", X"EA9", 
X"EA3", X"E9C", X"E94", X"E8D", X"E85", X"E7C", X"E73", X"E6A", 
X"E5F", X"E55", X"E4A", X"E3F", X"E33", X"E26", X"E19", X"E0C", 
X"DFF", X"DF0", X"DE1", X"DD2", X"DC3", X"DB3", X"DA2", X"D90", 
X"D80", X"D6E", X"D5B", X"D47", X"D35", X"D21", X"D0C", X"CF7", 
X"CE1", X"CCD", X"CB6", X"C9F", X"C87", X"C71", X"C59", X"C3F", 
X"C26", X"C0E", X"BF4", X"BD9", X"BBE", X"BA2", X"B88", X"B6B", 
X"B4E", X"B30", X"B15", X"AF7", X"AD8", X"AB8", X"A9B", X"A7B", 
X"A5B", X"A3A", X"A1B", X"9F9", X"9D7", X"9B5", X"992", X"971", 
X"94E", X"929", X"905", X"8E3", X"8BE", X"898", X"872", X"850", 
X"829", X"802", X"7DB", X"7B3", X"78F", X"766", X"73E", X"715", 
X"6EF", X"6C6", X"69C", X"672", X"64B", X"621", X"5F6", X"5CB", 
X"5A3", X"578", X"54C", X"520", X"4F4", X"4CB", X"49F", X"472", 
X"445", X"41C", X"3EE", X"3C1", X"393", X"369", X"33B", X"30D", 
X"2DF", X"2B0", X"286", X"257", X"229", X"1FA", X"1CF", X"1A0", 
X"171", X"142", X"117", X"0E8", X"0B9", X"089", X"05E", X"02F", 
X"000", X"FD0", X"FA1", X"F76", X"F46", X"F17", X"EE8", X"EBD", 
X"E8E", X"E5F", X"E30", X"E05", X"DD6", X"DA8", X"D79", X"D4F", 
X"D20", X"CF2", X"CC4", X"C96", X"C6C", X"C3E", X"C11", X"BE3", 
X"BBA", X"B8D", X"B60", X"B34", X"B0B", X"ADF", X"AB3", X"A87", 
X"A5C", X"A34", X"A09", X"9DE", X"9B4", X"98D", X"963", X"939", 
X"910", X"8EA", X"8C1", X"899", X"870", X"84C", X"824", X"7FD", 
X"7D6", X"7AF", X"78D", X"767", X"741", X"71C", X"6FA", X"6D6", 
X"6B1", X"68E", X"66D", X"64A", X"628", X"606", X"5E4", X"5C5", 
X"5A4", X"584", X"564", X"547", X"527", X"508", X"4EA", X"4CF", 
X"4B1", X"494", X"477", X"45D", X"441", X"426", X"40B", X"3F1", 
X"3D9", X"3C0", X"3A6", X"38E", X"378", X"360", X"349", X"332", 
X"31E", X"308", X"2F3", X"2DE", X"2CA", X"2B8", X"2A4", X"291", 
X"27F", X"26F", X"25D", X"24C", X"23C", X"22D", X"21E", X"20F", 
X"200", X"1F3", X"1E6", X"1D9", X"1CC", X"1C0", X"1B5", X"1AA", 
X"1A0", X"195", X"18C", X"183", X"17A", X"172", X"16B", X"163", 
X"15C", X"156", X"150", X"14B", X"146", X"141", X"13D", X"139", 
X"136", X"133", X"130", X"12E", X"12D", X"12C", X"12B", X"12A", 
X"12A", X"12B", X"12C", X"12D", X"12E", X"131", X"133", X"136", 
X"139", X"13C", X"140", X"145", X"149", X"14E", X"153", X"159", 
X"15F", X"165", X"16C", X"173", X"17A", X"181", X"189", X"192", 
X"19A", X"1A2", X"1AC", X"1B5", X"1BF", X"1C8", X"1D2", X"1DD", 
X"1E8", X"1F3", X"1FE", X"209", X"215", X"221", X"22C", X"239", 
X"246", X"253", X"25F", X"26C", X"27A", X"287", X"295", X"2A2", 
X"2B0", X"2BF", X"2CD", X"2DB", X"2EA", X"2F9", X"308", X"316", 
X"325", X"335", X"344", X"353", X"363", X"373", X"383", X"393", 
X"3A1", X"3B2", X"3C2", X"3D2", X"3E1", X"3F2", X"402", X"413", 
X"422", X"432", X"443", X"454", X"464", X"473", X"484", X"495", 
X"4A5", X"4B4", X"4C5", X"4D6", X"4E6", X"4F5", X"506", X"516", 
X"526", X"535", X"545", X"555", X"566", X"576", X"584", X"594", 
X"5A4", X"5B3", X"5C2", X"5D1", X"5E0", X"5F0", X"5FD", X"60C", 
X"61B", X"62A", X"639", X"646", X"655", X"663", X"671", X"67E", 
X"68C", X"699", X"6A7", X"6B3", X"6C0", X"6CD", X"6DA", X"6E6", 
X"6F2", X"6FF", X"70B", X"717", X"722", X"72E", X"739", X"744", 
X"74F", X"759", X"764", X"76F", X"778", X"783", X"78D", X"796", 
X"7A0", X"7A8", X"7B2", X"7BB", X"7C4", X"7CB", X"7D4", X"7DC", 
X"7E4", X"7EB", X"7F3", X"7FA", X"801", X"808", X"80E", X"815", 
X"81B", X"821", X"827", X"82D", X"832", X"837", X"83C", X"841", 
X"846", X"84A", X"84E", X"852", X"856", X"85A", X"85D", X"861", 
X"864", X"867", X"869", X"86C", X"86E", X"870", X"872", X"874", 
X"875", X"877", X"878", X"879", X"87A", X"87B", X"87B", X"87C", 
X"87C", X"87C", X"87C", X"87B", X"87B", X"87A", X"87A", X"879", 
X"878", X"876", X"875", X"874", X"872", X"870", X"86E", X"86C", 
X"86A", X"868", X"866", X"863", X"860", X"85E", X"85B", X"858", 
X"855", X"852", X"84E", X"84B", X"847", X"843", X"840", X"83C", 
X"838", X"834", X"831", X"82C", X"828", X"824", X"820", X"81B", 
X"817", X"812", X"80D", X"809", X"804", X"800", X"7FB", X"7F6", 
X"7F1", X"7EC", X"7E7", X"7E3", X"7DE", X"7D9", X"7D4", X"7CF", 
X"7CA", X"7C5", X"7BF", X"7BA", X"7B5", X"7B0", X"7AB", X"7A6", 
X"7A1", X"79C", X"797", X"791", X"78D", X"788", X"783", X"77D", 
X"778", X"774", X"76F", X"76A", X"765", X"760", X"75B", X"756", 
X"752", X"74D", X"749", X"744", X"73F", X"73B", X"737", X"732", 
X"72E", X"729", X"725", X"721", X"71D", X"719", X"715", X"711", 
X"70D", X"70A", X"706", X"703", X"6FF", X"6FB", X"6F8", X"6F5", 
X"6F2", X"6EE", X"6EB", X"6E9", X"6E6", X"6E3", X"6E0", X"6DD", 
X"6DB", X"6D8", X"6D6", X"6D4", X"6D2", X"6CF", X"6CD", X"6CB", 
X"6CA", X"6C8", X"6C6", X"6C5", X"6C3", X"6C2", X"6C1", X"6BF", 
X"6BE", X"6BD", X"6BD", X"6BC", X"6BB", X"6BA", X"6BA", X"6BA", 
X"6B9", X"6B9", X"6B9", X"6B9", X"6B9", X"6B9", X"6B9", X"6BA", 
X"6BA", X"6BB", X"6BB", X"6BC", X"6BD", X"6BE", X"6BE", X"6C0", 
X"6C1", X"6C2", X"6C3", X"6C5", X"6C6", X"6C8", X"6C9", X"6CB", 
X"6CD", X"6CF", X"6D1", X"6D3", X"6D5", X"6D7", X"6DA", X"6DC", 
X"6DE", X"6E1", X"6E4", X"6E6", X"6E9", X"6EC", X"6EF", X"6F2", 
X"6F5", X"6F8", X"6FB", X"6FE", X"701", X"705", X"708", X"70C", 
X"70F", X"713", X"716", X"71A", X"71E", X"722", X"726", X"72A", 
X"72E", X"731", X"736", X"73A", X"73E", X"742", X"746", X"74B", 
X"74F", X"753", X"758", X"75C", X"761", X"765", X"76A", X"76E", 
X"773", X"778", X"77C", X"781", X"786", X"78B", X"790", X"794", 
X"799", X"79F", X"7A3", X"7A8", X"7AD", X"7B2", X"7B7", X"7BC", 
X"7C1", X"7C7", X"7CC", X"7D1", X"7D6", X"7DB", X"7E1", X"7E5", 
X"7EB", X"7F0", X"7F6", X"7FA", X"800", X"805", X"80B", X"810", 
X"815", X"81B", X"820", X"826", X"82B", X"830", X"836", X"83B", 
X"840", X"846", X"84C", X"851", X"856", X"85C", X"862", X"867", 
X"86D", X"872", X"878", X"87D", X"883", X"888", X"88E", X"894", 
X"899", X"89F", X"8A4", X"8AA", X"8B0", X"8B6", X"8BB", X"8C1", 
X"8C7", X"8CC", X"8D2", X"8D8", X"8DD", X"8E3", X"8E9", X"8EF", 
X"8F5", X"8FB", X"900", X"906", X"90C", X"912", X"918", X"91E", 
X"924", X"92A", X"930", X"935", X"93C", X"942", X"948", X"94E", 
X"954", X"95A", X"960", X"967", X"96C", X"973", X"979", X"980", 
X"986", X"98C", X"993", X"999", X"99F", X"9A6", X"9AC", X"9B3", 
X"9B9", X"9C0", X"9C7", X"9CD", X"9D4", X"9DA", X"9E1", X"9E8", 
X"9EF", X"9F6", X"9FD", X"A04", X"A0B", X"A11", X"A19", X"A20", 
X"A27", X"A2E", X"A35", X"A3D", X"A44", X"A4C", X"A52", X"A5A", 
X"A62", X"A69", X"A70", X"A78", X"A80", X"A88", X"A8F", X"A97", 
X"A9F", X"AA7", X"AAF", X"AB6", X"ABE", X"AC6", X"ACF", X"AD6", 
X"ADF", X"AE7", X"AEF", X"AF7", X"B00", X"B08", X"B11", X"B19", 
X"B21", X"B2A", X"B33", X"B3C", X"B44", X"B4C", X"B55", X"B5E", 
X"B66", X"B70", X"B79", X"B82", X"B8A", X"B93", X"B9C", X"BA6", 
X"BAF", X"BB7", X"BC1", X"BCA", X"BD4", X"BDC", X"BE6", X"BEF", 
X"BF9", X"C01", X"C0B", X"C14", X"C1E", X"C28", X"C30", X"C3A", 
X"C44", X"C4D", X"C56", X"C60", X"C69", X"C73", X"C7C", X"C86", 
X"C8F", X"C99", X"CA2", X"CAC", X"CB5", X"CBF", X"CC9", X"CD2", 
X"CDB", X"CE5", X"CEF", X"CF7", X"D01", X"D0B", X"D14", X"D1D", 
X"D26", X"D30", X"D39", X"D43", X"D4B", X"D54", X"D5E", X"D67", 
X"D6F", X"D79", X"D82", X"D8B", X"D93", X"D9C", X"DA5", X"DAE", 
X"DB6", X"DBE", X"DC7", X"DD0", X"DD8", X"DE0", X"DE8", X"DF0", 
X"DF8", X"E00", X"E08", X"E10", X"E18", X"E1F", X"E26", X"E2E", 
X"E35", X"E3D", X"E43", X"E4A", X"E51", X"E58", X"E5E", X"E65", 
X"E6C", X"E72", X"E78", X"E7E", X"E84", X"E8A", X"E8F", X"E95", 
X"E9A", X"EA0", X"EA5", X"EAA", X"EAF", X"EB3", X"EB8", X"EBC", 
X"EC1", X"EC5", X"EC9", X"ECC", X"ED0", X"ED3", X"ED7", X"EDA", 
X"EDD", X"EE0", X"EE2", X"EE5", X"EE7", X"EE9", X"EEB", X"EED", 
X"EEE", X"EF0", X"EF1", X"EF2", X"EF3", X"EF3", X"EF4", X"EF4", 
X"EF4", X"EF4", X"EF4", X"EF3", X"EF2", X"EF2", X"EF0", X"EEF", 
X"EEE", X"EEC", X"EEA", X"EE8", X"EE6", X"EE3", X"EE0", X"EDD", 
X"EDA", X"ED7", X"ED4", X"ED0", X"ECC", X"EC8", X"EC4", X"EBF", 
X"EBA", X"EB5", X"EB0", X"EAB", X"EA5", X"E9F", X"E99", X"E93", 
X"E8D", X"E86", X"E7F", X"E79", X"E71", X"E6A", X"E62", X"E5B", 
X"E53", X"E4A", X"E42", X"E39", X"E31", X"E28", X"E1E", X"E15", 
X"E0C", X"E02", X"DF8", X"DEE", X"DE4", X"DDA", X"DCF", X"DC4", 
X"DBA", X"DAE", X"DA3", X"D97", X"D8B", X"D80", X"D74", X"D68", 
X"D5B", X"D50", X"D43", X"D36", X"D29", X"D1D", X"D0F", X"D02", 
X"CF4", X"CE6", X"CD9", X"CCB", X"CBD", X"CAF", X"CA1", X"C93", 
X"C84", X"C75", X"C68", X"C59", X"C49", X"C3A", X"C2C", X"C1D", 
X"C0D", X"BFE", X"BEE", X"BE0", X"BD0", X"BC0", X"BB0", X"BA1", 
X"B91", X"B81", X"B71", X"B62", X"B52", X"B41", X"B31", X"B21", 
X"B12", X"B01", X"AF1", X"AE0", X"AD1", X"AC1", X"AB0", X"AA0", 
X"A91", X"A80", X"A70", X"A5F", X"A50", X"A40", X"A2F", X"A1F", 
X"A0E", X"A00", X"9EF", X"9DF", X"9CF", X"9C0", X"9B0", X"9A0", 
X"990", X"982", X"972", X"963", X"953", X"943", X"935", X"926", 
X"917", X"908", X"8FA", X"8EB", X"8DC", X"8CE", X"8C0", X"8B2", 
X"8A4", X"896", X"889", X"87B", X"86D", X"860", X"852", X"846", 
X"839", X"82C", X"81F", X"814", X"808", X"7FB", X"7EF", X"7E4", 
X"7D9", X"7CD", X"7C2", X"7B7", X"7AD", X"7A2", X"798", X"78D", 
X"784", X"77A", X"771", X"767", X"75F", X"756", X"74D", X"744", 
X"73D", X"735", X"72D", X"725", X"71E", X"717", X"711", X"70A", 
X"704", X"6FE", X"6F8", X"6F2", X"6ED", X"6E8", X"6E3", X"6DF", 
X"6DA", X"6D6", X"6D3", X"6CF", X"6CC", X"6C9", X"6C6", X"6C4", 
X"6C1", X"6BF", X"6BE", X"6BC", X"6BB", X"6BA", X"6BA", X"6B9", 
X"6B9", X"6B9", X"6BA", X"6BA", X"6BB", X"6BC", X"6BE", X"6BF", 
X"6C1", X"6C4", X"6C6", X"6C9", X"6CC", X"6CF", X"6D3", X"6D6", 
X"6DA", X"6DF", X"6E3", X"6E8", X"6ED", X"6F2", X"6F8", X"6FE", 
X"704", X"70A", X"711", X"717", X"71E", X"725", X"72D", X"735", 
X"73D", X"744", X"74D", X"756", X"75F", X"767", X"771", X"77A", 
X"784", X"78D", X"798", X"7A2", X"7AD", X"7B7", X"7C2", X"7CD", 
X"7D9", X"7E4", X"7EF", X"7FB", X"808", X"814", X"81F", X"82C", 
X"839", X"846", X"852", X"860", X"86D", X"87B", X"889", X"896", 
X"8A4", X"8B2", X"8C0", X"8CE", X"8DC", X"8EB", X"8FA", X"908", 
X"917", X"926", X"935", X"943", X"953", X"963", X"972", X"982", 
X"990", X"9A0", X"9B0", X"9C0", X"9CF", X"9DF", X"9EF", X"A00", 
X"A0E", X"A1F", X"A2F", X"A40", X"A50", X"A5F", X"A70", X"A80", 
X"A91", X"AA0", X"AB0", X"AC1", X"AD1", X"AE0", X"AF1", X"B01", 
X"B12", X"B21", X"B31", X"B41", X"B52", X"B62", X"B71", X"B81", 
X"B91", X"BA1", X"BB0", X"BC0", X"BD0", X"BE0", X"BEE", X"BFE", 
X"C0D", X"C1D", X"C2C", X"C3A", X"C49", X"C59", X"C68", X"C75", 
X"C84", X"C93", X"CA1", X"CAF", X"CBD", X"CCB", X"CD9", X"CE6", 
X"CF4", X"D02", X"D0F", X"D1D", X"D29", X"D36", X"D43", X"D50", 
X"D5B", X"D68", X"D74", X"D80", X"D8B", X"D97", X"DA3", X"DAE", 
X"DBA", X"DC4", X"DCF", X"DDA", X"DE4", X"DEE", X"DF8", X"E02", 
X"E0C", X"E15", X"E1E", X"E28", X"E31", X"E39", X"E42", X"E4A", 
X"E53", X"E5B", X"E62", X"E6A", X"E71", X"E79", X"E7F", X"E86", 
X"E8D", X"E93", X"E99", X"E9F", X"EA5", X"EAB", X"EB0", X"EB5", 
X"EBA", X"EBF", X"EC4", X"EC8", X"ECC", X"ED0", X"ED4", X"ED7", 
X"EDA", X"EDD", X"EE0", X"EE3", X"EE6", X"EE8", X"EEA", X"EEC", 
X"EEE", X"EEF", X"EF0", X"EF2", X"EF2", X"EF3", X"EF4", X"EF4", 
X"EF4", X"EF4", X"EF4", X"EF3", X"EF3", X"EF2", X"EF1", X"EF0", 
X"EEE", X"EED", X"EEB", X"EE9", X"EE7", X"EE5", X"EE2", X"EE0", 
X"EDD", X"EDA", X"ED7", X"ED3", X"ED0", X"ECC", X"EC9", X"EC5", 
X"EC1", X"EBC", X"EB8", X"EB3", X"EAF", X"EAA", X"EA5", X"EA0", 
X"E9A", X"E95", X"E8F", X"E8A", X"E84", X"E7E", X"E78", X"E72", 
X"E6C", X"E65", X"E5E", X"E58", X"E51", X"E4A", X"E43", X"E3D", 
X"E35", X"E2E", X"E26", X"E1F", X"E18", X"E10", X"E08", X"E00", 
X"DF8", X"DF0", X"DE8", X"DE0", X"DD8", X"DD0", X"DC7", X"DBE", 
X"DB6", X"DAE", X"DA5", X"D9C", X"D93", X"D8B", X"D82", X"D79", 
X"D6F", X"D67", X"D5E", X"D54", X"D4B", X"D43", X"D39", X"D30", 
X"D26", X"D1D", X"D14", X"D0B", X"D01", X"CF7", X"CEF", X"CE5", 
X"CDB", X"CD2", X"CC9", X"CBF", X"CB5", X"CAC", X"CA2", X"C99", 
X"C8F", X"C86", X"C7C", X"C73", X"C69", X"C60", X"C56", X"C4D", 
X"C44", X"C3A", X"C30", X"C28", X"C1E", X"C14", X"C0B", X"C01", 
X"BF9", X"BEF", X"BE6", X"BDC", X"BD4", X"BCA", X"BC1", X"BB7", 
X"BAF", X"BA6", X"B9C", X"B93", X"B8A", X"B82", X"B79", X"B70", 
X"B66", X"B5E", X"B55", X"B4C", X"B44", X"B3C", X"B33", X"B2A", 
X"B21", X"B19", X"B11", X"B08", X"B00", X"AF7", X"AEF", X"AE7", 
X"ADF", X"AD6", X"ACF", X"AC6", X"ABE", X"AB6", X"AAF", X"AA7", 
X"A9F", X"A97", X"A8F", X"A88", X"A80", X"A78", X"A70", X"A69", 
X"A62", X"A5A", X"A52", X"A4C", X"A44", X"A3D", X"A35", X"A2E", 
X"A27", X"A20", X"A19", X"A11", X"A0B", X"A04", X"9FD", X"9F6", 
X"9EF", X"9E8", X"9E1", X"9DA", X"9D4", X"9CD", X"9C7", X"9C0", 
X"9B9", X"9B3", X"9AC", X"9A6", X"99F", X"999", X"993", X"98C", 
X"986", X"980", X"979", X"973", X"96C", X"967", X"960", X"95A", 
X"954", X"94E", X"948", X"942", X"93C", X"935", X"930", X"92A", 
X"924", X"91E", X"918", X"912", X"90C", X"906", X"900", X"8FB", 
X"8F5", X"8EF", X"8E9", X"8E3", X"8DD", X"8D8", X"8D2", X"8CC", 
X"8C7", X"8C1", X"8BB", X"8B6", X"8B0", X"8AA", X"8A4", X"89F", 
X"899", X"894", X"88E", X"888", X"883", X"87D", X"878", X"872", 
X"86D", X"867", X"862", X"85C", X"856", X"851", X"84C", X"846", 
X"840", X"83B", X"836", X"830", X"82B", X"826", X"820", X"81B", 
X"815", X"810", X"80B", X"805", X"800", X"7FA", X"7F6", X"7F0", 
X"7EB", X"7E5", X"7E1", X"7DB", X"7D6", X"7D1", X"7CC", X"7C7", 
X"7C1", X"7BC", X"7B7", X"7B2", X"7AD", X"7A8", X"7A3", X"79F", 
X"799", X"794", X"790", X"78B", X"786", X"781", X"77C", X"778", 
X"773", X"76E", X"76A", X"765", X"761", X"75C", X"758", X"753", 
X"74F", X"74B", X"746", X"742", X"73E", X"73A", X"736", X"731", 
X"72D", X"72A", X"726", X"722", X"71E", X"71A", X"716", X"713", 
X"70F", X"70C", X"708", X"705", X"701", X"6FE", X"6FB", X"6F8", 
X"6F5", X"6F2", X"6EF", X"6EC", X"6E9", X"6E6", X"6E4", X"6E1", 
X"6DE", X"6DC", X"6DA", X"6D7", X"6D5", X"6D3", X"6D1", X"6CF", 
X"6CD", X"6CB", X"6C9", X"6C8", X"6C6", X"6C5", X"6C3", X"6C2", 
X"6C1", X"6C0", X"6BE", X"6BE", X"6BD", X"6BC", X"6BB", X"6BB", 
X"6BA", X"6BA", X"6B9", X"6B9", X"6B9", X"6B9", X"6B9", X"6B9", 
X"6B9", X"6BA", X"6BA", X"6BA", X"6BB", X"6BC", X"6BD", X"6BD", 
X"6BE", X"6BF", X"6C1", X"6C2", X"6C3", X"6C5", X"6C6", X"6C8", 
X"6CA", X"6CB", X"6CD", X"6CF", X"6D2", X"6D4", X"6D6", X"6D8", 
X"6DB", X"6DD", X"6E0", X"6E3", X"6E6", X"6E9", X"6EB", X"6EE", 
X"6F2", X"6F5", X"6F8", X"6FB", X"6FF", X"703", X"706", X"70A", 
X"70D", X"711", X"715", X"719", X"71D", X"721", X"725", X"729", 
X"72E", X"732", X"737", X"73B", X"73F", X"744", X"749", X"74D", 
X"752", X"756", X"75B", X"760", X"765", X"76A", X"76F", X"774", 
X"778", X"77D", X"783", X"788", X"78D", X"791", X"797", X"79C", 
X"7A1", X"7A6", X"7AB", X"7B0", X"7B5", X"7BA", X"7BF", X"7C5", 
X"7CA", X"7CF", X"7D4", X"7D9", X"7DE", X"7E3", X"7E7", X"7EC", 
X"7F1", X"7F6", X"7FB", X"800", X"804", X"809", X"80D", X"812", 
X"817", X"81B", X"820", X"824", X"828", X"82C", X"831", X"834", 
X"838", X"83C", X"840", X"843", X"847", X"84B", X"84E", X"852", 
X"855", X"858", X"85B", X"85E", X"860", X"863", X"866", X"868", 
X"86A", X"86C", X"86E", X"870", X"872", X"874", X"875", X"876", 
X"878", X"879", X"87A", X"87A", X"87B", X"87B", X"87C", X"87C", 
X"87C", X"87C", X"87B", X"87B", X"87A", X"879", X"878", X"877", 
X"875", X"874", X"872", X"870", X"86E", X"86C", X"869", X"867", 
X"864", X"861", X"85D", X"85A", X"856", X"852", X"84E", X"84A", 
X"846", X"841", X"83C", X"837", X"832", X"82D", X"827", X"821", 
X"81B", X"815", X"80E", X"808", X"801", X"7FA", X"7F3", X"7EB", 
X"7E4", X"7DC", X"7D4", X"7CB", X"7C4", X"7BB", X"7B2", X"7A8", 
X"7A0", X"796", X"78D", X"783", X"778", X"76F", X"764", X"759", 
X"74F", X"744", X"739", X"72E", X"722", X"717", X"70B", X"6FF", 
X"6F2", X"6E6", X"6DA", X"6CD", X"6C0", X"6B3", X"6A7", X"699", 
X"68C", X"67E", X"671", X"663", X"655", X"646", X"639", X"62A", 
X"61B", X"60C", X"5FD", X"5F0", X"5E0", X"5D1", X"5C2", X"5B3", 
X"5A4", X"594", X"584", X"576", X"566", X"555", X"545", X"535", 
X"526", X"516", X"506", X"4F5", X"4E6", X"4D6", X"4C5", X"4B4", 
X"4A5", X"495", X"484", X"473", X"464", X"454", X"443", X"432", 
X"422", X"413", X"402", X"3F2", X"3E1", X"3D2", X"3C2", X"3B2", 
X"3A1", X"393", X"383", X"373", X"363", X"353", X"344", X"335", 
X"325", X"316", X"308", X"2F9", X"2EA", X"2DB", X"2CD", X"2BF", 
X"2B0", X"2A2", X"295", X"287", X"27A", X"26C", X"25F", X"253", 
X"246", X"239", X"22C", X"221", X"215", X"209", X"1FE", X"1F3", 
X"1E8", X"1DD", X"1D2", X"1C8", X"1BF", X"1B5", X"1AC", X"1A2", 
X"19A", X"192", X"189", X"181", X"17A", X"173", X"16C", X"165", 
X"15F", X"159", X"153", X"14E", X"149", X"145", X"140", X"13C", 
X"139", X"136", X"133", X"131", X"12E", X"12D", X"12C", X"12B", 
X"12A", X"12A", X"12B", X"12C", X"12D", X"12E", X"130", X"133", 
X"136", X"139", X"13D", X"141", X"146", X"14B", X"150", X"156", 
X"15C", X"163", X"16B", X"172", X"17A", X"183", X"18C", X"195", 
X"1A0", X"1AA", X"1B5", X"1C0", X"1CC", X"1D9", X"1E6", X"1F3", 
X"200", X"20F", X"21E", X"22D", X"23C", X"24C", X"25D", X"26F", 
X"27F", X"291", X"2A4", X"2B8", X"2CA", X"2DE", X"2F3", X"308", 
X"31E", X"332", X"349", X"360", X"378", X"38E", X"3A6", X"3C0", 
X"3D9", X"3F1", X"40B", X"426", X"441", X"45D", X"477", X"494", 
X"4B1", X"4CF", X"4EA", X"508", X"527", X"547", X"564", X"584", 
X"5A4", X"5C5", X"5E4", X"606", X"628", X"64A", X"66D", X"68E", 
X"6B1", X"6D6", X"6FA", X"71C", X"741", X"767", X"78D", X"7AF", 
X"7D6", X"7FD", X"824", X"84C", X"870", X"899", X"8C1", X"8EA", 
X"910", X"939", X"963", X"98D", X"9B4", X"9DE", X"A09", X"A34", 
X"A5C", X"A87", X"AB3", X"ADF", X"B0B", X"B34", X"B60", X"B8D", 
X"BBA", X"BE3", X"C11", X"C3E", X"C6C", X"C96", X"CC4", X"CF2", 
X"D20", X"D4F", X"D79", X"DA8", X"DD6", X"E05", X"E30", X"E5F", 
X"E8E", X"EBD", X"EE8", X"F17", X"F46", X"F76", X"FA1", X"FD0"
);

signal data : std_logic_vector(31 downto 0);
signal unsignedIndex : unsigned(11 downto 0) := X"000";

begin

rom_select: process (clk, en)
begin
	if (rising_edge(clk)) then
    if (en = '1') then
		unsignedIndex <= unsigned(address_reg);
		data <= (SIN_ROM(to_integer(unsignedIndex)) & x"00000");
		sin_out <= std_logic_vector(shift_right(signed(data), 20));
    end if;
  end if;
end process rom_select;

end rtl;
