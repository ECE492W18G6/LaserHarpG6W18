-- soc_system.vhd

-- Generated using ACDS version 17.0 602

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity soc_system is
	port (
		audio_0_external_interface_ADCDAT                : in    std_logic                     := '0';             --                  audio_0_external_interface.ADCDAT
		audio_0_external_interface_ADCLRCK               : in    std_logic                     := '0';             --                                            .ADCLRCK
		audio_0_external_interface_BCLK                  : in    std_logic                     := '0';             --                                            .BCLK
		audio_0_external_interface_DACDAT                : out   std_logic;                                        --                                            .DACDAT
		audio_0_external_interface_DACLRCK               : in    std_logic                     := '0';             --                                            .DACLRCK
		audio_and_video_config_0_external_interface_SDAT : inout std_logic                     := '0';             -- audio_and_video_config_0_external_interface.SDAT
		audio_and_video_config_0_external_interface_SCLK : out   std_logic;                                        --                                            .SCLK
		buttons_external_connection_export               : in    std_logic_vector(3 downto 0)  := (others => '0'); --                 buttons_external_connection.export
		character_lcd_0_external_interface_DATA          : inout std_logic_vector(7 downto 0)  := (others => '0'); --          character_lcd_0_external_interface.DATA
		character_lcd_0_external_interface_ON            : out   std_logic;                                        --                                            .ON
		character_lcd_0_external_interface_BLON          : out   std_logic;                                        --                                            .BLON
		character_lcd_0_external_interface_EN            : out   std_logic;                                        --                                            .EN
		character_lcd_0_external_interface_RS            : out   std_logic;                                        --                                            .RS
		character_lcd_0_external_interface_RW            : out   std_logic;                                        --                                            .RW
		clk_clk                                          : in    std_logic                     := '0';             --                                         clk.clk
		hps_io_hps_io_emac1_inst_TX_CLK                  : out   std_logic;                                        --                                      hps_io.hps_io_emac1_inst_TX_CLK
		hps_io_hps_io_emac1_inst_TXD0                    : out   std_logic;                                        --                                            .hps_io_emac1_inst_TXD0
		hps_io_hps_io_emac1_inst_TXD1                    : out   std_logic;                                        --                                            .hps_io_emac1_inst_TXD1
		hps_io_hps_io_emac1_inst_TXD2                    : out   std_logic;                                        --                                            .hps_io_emac1_inst_TXD2
		hps_io_hps_io_emac1_inst_TXD3                    : out   std_logic;                                        --                                            .hps_io_emac1_inst_TXD3
		hps_io_hps_io_emac1_inst_RXD0                    : in    std_logic                     := '0';             --                                            .hps_io_emac1_inst_RXD0
		hps_io_hps_io_emac1_inst_MDIO                    : inout std_logic                     := '0';             --                                            .hps_io_emac1_inst_MDIO
		hps_io_hps_io_emac1_inst_MDC                     : out   std_logic;                                        --                                            .hps_io_emac1_inst_MDC
		hps_io_hps_io_emac1_inst_RX_CTL                  : in    std_logic                     := '0';             --                                            .hps_io_emac1_inst_RX_CTL
		hps_io_hps_io_emac1_inst_TX_CTL                  : out   std_logic;                                        --                                            .hps_io_emac1_inst_TX_CTL
		hps_io_hps_io_emac1_inst_RX_CLK                  : in    std_logic                     := '0';             --                                            .hps_io_emac1_inst_RX_CLK
		hps_io_hps_io_emac1_inst_RXD1                    : in    std_logic                     := '0';             --                                            .hps_io_emac1_inst_RXD1
		hps_io_hps_io_emac1_inst_RXD2                    : in    std_logic                     := '0';             --                                            .hps_io_emac1_inst_RXD2
		hps_io_hps_io_emac1_inst_RXD3                    : in    std_logic                     := '0';             --                                            .hps_io_emac1_inst_RXD3
		hps_io_hps_io_sdio_inst_CMD                      : inout std_logic                     := '0';             --                                            .hps_io_sdio_inst_CMD
		hps_io_hps_io_sdio_inst_D0                       : inout std_logic                     := '0';             --                                            .hps_io_sdio_inst_D0
		hps_io_hps_io_sdio_inst_D1                       : inout std_logic                     := '0';             --                                            .hps_io_sdio_inst_D1
		hps_io_hps_io_sdio_inst_CLK                      : out   std_logic;                                        --                                            .hps_io_sdio_inst_CLK
		hps_io_hps_io_sdio_inst_D2                       : inout std_logic                     := '0';             --                                            .hps_io_sdio_inst_D2
		hps_io_hps_io_sdio_inst_D3                       : inout std_logic                     := '0';             --                                            .hps_io_sdio_inst_D3
		hps_io_hps_io_usb1_inst_D0                       : inout std_logic                     := '0';             --                                            .hps_io_usb1_inst_D0
		hps_io_hps_io_usb1_inst_D1                       : inout std_logic                     := '0';             --                                            .hps_io_usb1_inst_D1
		hps_io_hps_io_usb1_inst_D2                       : inout std_logic                     := '0';             --                                            .hps_io_usb1_inst_D2
		hps_io_hps_io_usb1_inst_D3                       : inout std_logic                     := '0';             --                                            .hps_io_usb1_inst_D3
		hps_io_hps_io_usb1_inst_D4                       : inout std_logic                     := '0';             --                                            .hps_io_usb1_inst_D4
		hps_io_hps_io_usb1_inst_D5                       : inout std_logic                     := '0';             --                                            .hps_io_usb1_inst_D5
		hps_io_hps_io_usb1_inst_D6                       : inout std_logic                     := '0';             --                                            .hps_io_usb1_inst_D6
		hps_io_hps_io_usb1_inst_D7                       : inout std_logic                     := '0';             --                                            .hps_io_usb1_inst_D7
		hps_io_hps_io_usb1_inst_CLK                      : in    std_logic                     := '0';             --                                            .hps_io_usb1_inst_CLK
		hps_io_hps_io_usb1_inst_STP                      : out   std_logic;                                        --                                            .hps_io_usb1_inst_STP
		hps_io_hps_io_usb1_inst_DIR                      : in    std_logic                     := '0';             --                                            .hps_io_usb1_inst_DIR
		hps_io_hps_io_usb1_inst_NXT                      : in    std_logic                     := '0';             --                                            .hps_io_usb1_inst_NXT
		hps_io_hps_io_spim1_inst_CLK                     : out   std_logic;                                        --                                            .hps_io_spim1_inst_CLK
		hps_io_hps_io_spim1_inst_MOSI                    : out   std_logic;                                        --                                            .hps_io_spim1_inst_MOSI
		hps_io_hps_io_spim1_inst_MISO                    : in    std_logic                     := '0';             --                                            .hps_io_spim1_inst_MISO
		hps_io_hps_io_spim1_inst_SS0                     : out   std_logic;                                        --                                            .hps_io_spim1_inst_SS0
		hps_io_hps_io_uart0_inst_RX                      : in    std_logic                     := '0';             --                                            .hps_io_uart0_inst_RX
		hps_io_hps_io_uart0_inst_TX                      : out   std_logic;                                        --                                            .hps_io_uart0_inst_TX
		hps_io_hps_io_i2c0_inst_SDA                      : inout std_logic                     := '0';             --                                            .hps_io_i2c0_inst_SDA
		hps_io_hps_io_i2c0_inst_SCL                      : inout std_logic                     := '0';             --                                            .hps_io_i2c0_inst_SCL
		hps_io_hps_io_i2c1_inst_SDA                      : inout std_logic                     := '0';             --                                            .hps_io_i2c1_inst_SDA
		hps_io_hps_io_i2c1_inst_SCL                      : inout std_logic                     := '0';             --                                            .hps_io_i2c1_inst_SCL
		hps_io_hps_io_gpio_inst_GPIO09                   : inout std_logic                     := '0';             --                                            .hps_io_gpio_inst_GPIO09
		hps_io_hps_io_gpio_inst_GPIO35                   : inout std_logic                     := '0';             --                                            .hps_io_gpio_inst_GPIO35
		hps_io_hps_io_gpio_inst_GPIO40                   : inout std_logic                     := '0';             --                                            .hps_io_gpio_inst_GPIO40
		hps_io_hps_io_gpio_inst_GPIO48                   : inout std_logic                     := '0';             --                                            .hps_io_gpio_inst_GPIO48
		hps_io_hps_io_gpio_inst_GPIO53                   : inout std_logic                     := '0';             --                                            .hps_io_gpio_inst_GPIO53
		hps_io_hps_io_gpio_inst_GPIO54                   : inout std_logic                     := '0';             --                                            .hps_io_gpio_inst_GPIO54
		hps_io_hps_io_gpio_inst_GPIO61                   : inout std_logic                     := '0';             --                                            .hps_io_gpio_inst_GPIO61
		memory_mem_a                                     : out   std_logic_vector(14 downto 0);                    --                                      memory.mem_a
		memory_mem_ba                                    : out   std_logic_vector(2 downto 0);                     --                                            .mem_ba
		memory_mem_ck                                    : out   std_logic;                                        --                                            .mem_ck
		memory_mem_ck_n                                  : out   std_logic;                                        --                                            .mem_ck_n
		memory_mem_cke                                   : out   std_logic;                                        --                                            .mem_cke
		memory_mem_cs_n                                  : out   std_logic;                                        --                                            .mem_cs_n
		memory_mem_ras_n                                 : out   std_logic;                                        --                                            .mem_ras_n
		memory_mem_cas_n                                 : out   std_logic;                                        --                                            .mem_cas_n
		memory_mem_we_n                                  : out   std_logic;                                        --                                            .mem_we_n
		memory_mem_reset_n                               : out   std_logic;                                        --                                            .mem_reset_n
		memory_mem_dq                                    : inout std_logic_vector(31 downto 0) := (others => '0'); --                                            .mem_dq
		memory_mem_dqs                                   : inout std_logic_vector(3 downto 0)  := (others => '0'); --                                            .mem_dqs
		memory_mem_dqs_n                                 : inout std_logic_vector(3 downto 0)  := (others => '0'); --                                            .mem_dqs_n
		memory_mem_odt                                   : out   std_logic;                                        --                                            .mem_odt
		memory_mem_dm                                    : out   std_logic_vector(3 downto 0);                     --                                            .mem_dm
		memory_oct_rzqin                                 : in    std_logic                     := '0';             --                                            .oct_rzqin
		photodiode_0_conduit_end_export0                 : in    std_logic                     := '0';             --                    photodiode_0_conduit_end.export0
		photodiode_0_conduit_end_export1                 : in    std_logic                     := '0';             --                                            .export1
		photodiode_0_conduit_end_export2                 : in    std_logic                     := '0';             --                                            .export2
		photodiode_0_conduit_end_export3                 : in    std_logic                     := '0';             --                                            .export3
		photodiode_0_conduit_end_export4                 : in    std_logic                     := '0';             --                                            .export4
		photodiode_0_conduit_end_export5                 : in    std_logic                     := '0';             --                                            .export5
		photodiode_0_conduit_end_export6                 : in    std_logic                     := '0';             --                                            .export6
		photodiode_0_conduit_end_export7                 : in    std_logic                     := '0';             --                                            .export7
		pll_0_outclk0_clk                                : out   std_logic;                                        --                               pll_0_outclk0.clk
		red_leds_external_connection_export              : out   std_logic_vector(9 downto 0);                     --                red_leds_external_connection.export
		reset_reset_n                                    : in    std_logic                     := '0';             --                                       reset.reset_n
		switches_external_connection_export              : in    std_logic_vector(9 downto 0)  := (others => '0')  --                switches_external_connection.export
	);
end entity soc_system;

architecture rtl of soc_system is
	component EnvelopeController is
		port (
			data_out : out std_logic_vector(31 downto 0);                    -- readdata
			read     : in  std_logic                     := 'X';             -- read
			write    : in  std_logic                     := 'X';             -- write
			data_in  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			reset    : in  std_logic                     := 'X';             -- reset
			clk      : in  std_logic                     := 'X'              -- clk
		);
	end component EnvelopeController;

	component synthesizer is
		port (
			clk       : in  std_logic                     := 'X';             -- clk
			reset     : in  std_logic                     := 'X';             -- reset
			phase_reg : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			data_out  : out std_logic_vector(31 downto 0);                    -- readdata
			read      : in  std_logic                     := 'X';             -- read
			write     : in  std_logic                     := 'X'              -- write
		);
	end component synthesizer;

	component soc_system_audio_0 is
		port (
			clk         : in  std_logic                     := 'X';             -- clk
			reset       : in  std_logic                     := 'X';             -- reset
			address     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			chipselect  : in  std_logic                     := 'X';             -- chipselect
			read        : in  std_logic                     := 'X';             -- read
			write       : in  std_logic                     := 'X';             -- write
			writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			irq         : out std_logic;                                        -- irq
			AUD_ADCDAT  : in  std_logic                     := 'X';             -- export
			AUD_ADCLRCK : in  std_logic                     := 'X';             -- export
			AUD_BCLK    : in  std_logic                     := 'X';             -- export
			AUD_DACDAT  : out std_logic;                                        -- export
			AUD_DACLRCK : in  std_logic                     := 'X'              -- export
		);
	end component soc_system_audio_0;

	component soc_system_audio_and_video_config_0 is
		port (
			clk         : in    std_logic                     := 'X';             -- clk
			reset       : in    std_logic                     := 'X';             -- reset
			address     : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			byteenable  : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			read        : in    std_logic                     := 'X';             -- read
			write       : in    std_logic                     := 'X';             -- write
			writedata   : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata    : out   std_logic_vector(31 downto 0);                    -- readdata
			waitrequest : out   std_logic;                                        -- waitrequest
			I2C_SDAT    : inout std_logic                     := 'X';             -- export
			I2C_SCLK    : out   std_logic                                         -- export
		);
	end component soc_system_audio_and_video_config_0;

	component soc_system_buttons is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- export
			irq        : out std_logic                                         -- irq
		);
	end component soc_system_buttons;

	component soc_system_character_lcd_0 is
		port (
			clk         : in    std_logic                    := 'X';             -- clk
			reset       : in    std_logic                    := 'X';             -- reset
			address     : in    std_logic                    := 'X';             -- address
			chipselect  : in    std_logic                    := 'X';             -- chipselect
			read        : in    std_logic                    := 'X';             -- read
			write       : in    std_logic                    := 'X';             -- write
			writedata   : in    std_logic_vector(7 downto 0) := (others => 'X'); -- writedata
			readdata    : out   std_logic_vector(7 downto 0);                    -- readdata
			waitrequest : out   std_logic;                                       -- waitrequest
			LCD_DATA    : inout std_logic_vector(7 downto 0) := (others => 'X'); -- export
			LCD_ON      : out   std_logic;                                       -- export
			LCD_BLON    : out   std_logic;                                       -- export
			LCD_EN      : out   std_logic;                                       -- export
			LCD_RS      : out   std_logic;                                       -- export
			LCD_RW      : out   std_logic                                        -- export
		);
	end component soc_system_character_lcd_0;

	component soc_system_hps_0 is
		generic (
			F2S_Width : integer := 2;
			S2F_Width : integer := 2
		);
		port (
			mem_a                    : out   std_logic_vector(14 downto 0);                    -- mem_a
			mem_ba                   : out   std_logic_vector(2 downto 0);                     -- mem_ba
			mem_ck                   : out   std_logic;                                        -- mem_ck
			mem_ck_n                 : out   std_logic;                                        -- mem_ck_n
			mem_cke                  : out   std_logic;                                        -- mem_cke
			mem_cs_n                 : out   std_logic;                                        -- mem_cs_n
			mem_ras_n                : out   std_logic;                                        -- mem_ras_n
			mem_cas_n                : out   std_logic;                                        -- mem_cas_n
			mem_we_n                 : out   std_logic;                                        -- mem_we_n
			mem_reset_n              : out   std_logic;                                        -- mem_reset_n
			mem_dq                   : inout std_logic_vector(31 downto 0) := (others => 'X'); -- mem_dq
			mem_dqs                  : inout std_logic_vector(3 downto 0)  := (others => 'X'); -- mem_dqs
			mem_dqs_n                : inout std_logic_vector(3 downto 0)  := (others => 'X'); -- mem_dqs_n
			mem_odt                  : out   std_logic;                                        -- mem_odt
			mem_dm                   : out   std_logic_vector(3 downto 0);                     -- mem_dm
			oct_rzqin                : in    std_logic                     := 'X';             -- oct_rzqin
			hps_io_emac1_inst_TX_CLK : out   std_logic;                                        -- hps_io_emac1_inst_TX_CLK
			hps_io_emac1_inst_TXD0   : out   std_logic;                                        -- hps_io_emac1_inst_TXD0
			hps_io_emac1_inst_TXD1   : out   std_logic;                                        -- hps_io_emac1_inst_TXD1
			hps_io_emac1_inst_TXD2   : out   std_logic;                                        -- hps_io_emac1_inst_TXD2
			hps_io_emac1_inst_TXD3   : out   std_logic;                                        -- hps_io_emac1_inst_TXD3
			hps_io_emac1_inst_RXD0   : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RXD0
			hps_io_emac1_inst_MDIO   : inout std_logic                     := 'X';             -- hps_io_emac1_inst_MDIO
			hps_io_emac1_inst_MDC    : out   std_logic;                                        -- hps_io_emac1_inst_MDC
			hps_io_emac1_inst_RX_CTL : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RX_CTL
			hps_io_emac1_inst_TX_CTL : out   std_logic;                                        -- hps_io_emac1_inst_TX_CTL
			hps_io_emac1_inst_RX_CLK : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RX_CLK
			hps_io_emac1_inst_RXD1   : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RXD1
			hps_io_emac1_inst_RXD2   : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RXD2
			hps_io_emac1_inst_RXD3   : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RXD3
			hps_io_sdio_inst_CMD     : inout std_logic                     := 'X';             -- hps_io_sdio_inst_CMD
			hps_io_sdio_inst_D0      : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D0
			hps_io_sdio_inst_D1      : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D1
			hps_io_sdio_inst_CLK     : out   std_logic;                                        -- hps_io_sdio_inst_CLK
			hps_io_sdio_inst_D2      : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D2
			hps_io_sdio_inst_D3      : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D3
			hps_io_usb1_inst_D0      : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D0
			hps_io_usb1_inst_D1      : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D1
			hps_io_usb1_inst_D2      : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D2
			hps_io_usb1_inst_D3      : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D3
			hps_io_usb1_inst_D4      : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D4
			hps_io_usb1_inst_D5      : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D5
			hps_io_usb1_inst_D6      : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D6
			hps_io_usb1_inst_D7      : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D7
			hps_io_usb1_inst_CLK     : in    std_logic                     := 'X';             -- hps_io_usb1_inst_CLK
			hps_io_usb1_inst_STP     : out   std_logic;                                        -- hps_io_usb1_inst_STP
			hps_io_usb1_inst_DIR     : in    std_logic                     := 'X';             -- hps_io_usb1_inst_DIR
			hps_io_usb1_inst_NXT     : in    std_logic                     := 'X';             -- hps_io_usb1_inst_NXT
			hps_io_spim1_inst_CLK    : out   std_logic;                                        -- hps_io_spim1_inst_CLK
			hps_io_spim1_inst_MOSI   : out   std_logic;                                        -- hps_io_spim1_inst_MOSI
			hps_io_spim1_inst_MISO   : in    std_logic                     := 'X';             -- hps_io_spim1_inst_MISO
			hps_io_spim1_inst_SS0    : out   std_logic;                                        -- hps_io_spim1_inst_SS0
			hps_io_uart0_inst_RX     : in    std_logic                     := 'X';             -- hps_io_uart0_inst_RX
			hps_io_uart0_inst_TX     : out   std_logic;                                        -- hps_io_uart0_inst_TX
			hps_io_i2c0_inst_SDA     : inout std_logic                     := 'X';             -- hps_io_i2c0_inst_SDA
			hps_io_i2c0_inst_SCL     : inout std_logic                     := 'X';             -- hps_io_i2c0_inst_SCL
			hps_io_i2c1_inst_SDA     : inout std_logic                     := 'X';             -- hps_io_i2c1_inst_SDA
			hps_io_i2c1_inst_SCL     : inout std_logic                     := 'X';             -- hps_io_i2c1_inst_SCL
			hps_io_gpio_inst_GPIO09  : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO09
			hps_io_gpio_inst_GPIO35  : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO35
			hps_io_gpio_inst_GPIO40  : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO40
			hps_io_gpio_inst_GPIO48  : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO48
			hps_io_gpio_inst_GPIO53  : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO53
			hps_io_gpio_inst_GPIO54  : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO54
			hps_io_gpio_inst_GPIO61  : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO61
			h2f_rst_n                : out   std_logic;                                        -- reset_n
			h2f_lw_axi_clk           : in    std_logic                     := 'X';             -- clk
			h2f_lw_AWID              : out   std_logic_vector(11 downto 0);                    -- awid
			h2f_lw_AWADDR            : out   std_logic_vector(20 downto 0);                    -- awaddr
			h2f_lw_AWLEN             : out   std_logic_vector(3 downto 0);                     -- awlen
			h2f_lw_AWSIZE            : out   std_logic_vector(2 downto 0);                     -- awsize
			h2f_lw_AWBURST           : out   std_logic_vector(1 downto 0);                     -- awburst
			h2f_lw_AWLOCK            : out   std_logic_vector(1 downto 0);                     -- awlock
			h2f_lw_AWCACHE           : out   std_logic_vector(3 downto 0);                     -- awcache
			h2f_lw_AWPROT            : out   std_logic_vector(2 downto 0);                     -- awprot
			h2f_lw_AWVALID           : out   std_logic;                                        -- awvalid
			h2f_lw_AWREADY           : in    std_logic                     := 'X';             -- awready
			h2f_lw_WID               : out   std_logic_vector(11 downto 0);                    -- wid
			h2f_lw_WDATA             : out   std_logic_vector(31 downto 0);                    -- wdata
			h2f_lw_WSTRB             : out   std_logic_vector(3 downto 0);                     -- wstrb
			h2f_lw_WLAST             : out   std_logic;                                        -- wlast
			h2f_lw_WVALID            : out   std_logic;                                        -- wvalid
			h2f_lw_WREADY            : in    std_logic                     := 'X';             -- wready
			h2f_lw_BID               : in    std_logic_vector(11 downto 0) := (others => 'X'); -- bid
			h2f_lw_BRESP             : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- bresp
			h2f_lw_BVALID            : in    std_logic                     := 'X';             -- bvalid
			h2f_lw_BREADY            : out   std_logic;                                        -- bready
			h2f_lw_ARID              : out   std_logic_vector(11 downto 0);                    -- arid
			h2f_lw_ARADDR            : out   std_logic_vector(20 downto 0);                    -- araddr
			h2f_lw_ARLEN             : out   std_logic_vector(3 downto 0);                     -- arlen
			h2f_lw_ARSIZE            : out   std_logic_vector(2 downto 0);                     -- arsize
			h2f_lw_ARBURST           : out   std_logic_vector(1 downto 0);                     -- arburst
			h2f_lw_ARLOCK            : out   std_logic_vector(1 downto 0);                     -- arlock
			h2f_lw_ARCACHE           : out   std_logic_vector(3 downto 0);                     -- arcache
			h2f_lw_ARPROT            : out   std_logic_vector(2 downto 0);                     -- arprot
			h2f_lw_ARVALID           : out   std_logic;                                        -- arvalid
			h2f_lw_ARREADY           : in    std_logic                     := 'X';             -- arready
			h2f_lw_RID               : in    std_logic_vector(11 downto 0) := (others => 'X'); -- rid
			h2f_lw_RDATA             : in    std_logic_vector(31 downto 0) := (others => 'X'); -- rdata
			h2f_lw_RRESP             : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- rresp
			h2f_lw_RLAST             : in    std_logic                     := 'X';             -- rlast
			h2f_lw_RVALID            : in    std_logic                     := 'X';             -- rvalid
			h2f_lw_RREADY            : out   std_logic;                                        -- rready
			f2h_irq_p0               : in    std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			f2h_irq_p1               : in    std_logic_vector(31 downto 0) := (others => 'X')  -- irq
		);
	end component soc_system_hps_0;

	component photodiode is
		port (
			avalon_slave_readdata : out std_logic_vector(7 downto 0);        -- readdata
			avalon_slave_read_n   : in  std_logic                    := 'X'; -- read_n
			conduit_end_0         : in  std_logic                    := 'X'; -- export0
			conduit_end_1         : in  std_logic                    := 'X'; -- export1
			conduit_end_2         : in  std_logic                    := 'X'; -- export2
			conduit_end_3         : in  std_logic                    := 'X'; -- export3
			conduit_end_4         : in  std_logic                    := 'X'; -- export4
			conduit_end_5         : in  std_logic                    := 'X'; -- export5
			conduit_end_6         : in  std_logic                    := 'X'; -- export6
			conduit_end_7         : in  std_logic                    := 'X'; -- export7
			clk                   : in  std_logic                    := 'X'; -- clk
			reset_n               : in  std_logic                    := 'X'  -- reset_n
		);
	end component photodiode;

	component soc_system_pll_0 is
		port (
			refclk   : in  std_logic := 'X'; -- clk
			rst      : in  std_logic := 'X'; -- reset
			outclk_0 : out std_logic;        -- clk
			locked   : out std_logic         -- export
		);
	end component soc_system_pll_0;

	component soc_system_red_leds is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(9 downto 0)                      -- export
		);
	end component soc_system_red_leds;

	component soc_system_switches is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- export
			irq        : out std_logic                                         -- irq
		);
	end component soc_system_switches;

	component soc_system_sysid_qsys_0 is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component soc_system_sysid_qsys_0;

	component soc_system_mm_interconnect_0 is
		port (
			hps_0_h2f_lw_axi_master_awid                                        : in  std_logic_vector(11 downto 0) := (others => 'X'); -- awid
			hps_0_h2f_lw_axi_master_awaddr                                      : in  std_logic_vector(20 downto 0) := (others => 'X'); -- awaddr
			hps_0_h2f_lw_axi_master_awlen                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awlen
			hps_0_h2f_lw_axi_master_awsize                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awsize
			hps_0_h2f_lw_axi_master_awburst                                     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- awburst
			hps_0_h2f_lw_axi_master_awlock                                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- awlock
			hps_0_h2f_lw_axi_master_awcache                                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awcache
			hps_0_h2f_lw_axi_master_awprot                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awprot
			hps_0_h2f_lw_axi_master_awvalid                                     : in  std_logic                     := 'X';             -- awvalid
			hps_0_h2f_lw_axi_master_awready                                     : out std_logic;                                        -- awready
			hps_0_h2f_lw_axi_master_wid                                         : in  std_logic_vector(11 downto 0) := (others => 'X'); -- wid
			hps_0_h2f_lw_axi_master_wdata                                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wdata
			hps_0_h2f_lw_axi_master_wstrb                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- wstrb
			hps_0_h2f_lw_axi_master_wlast                                       : in  std_logic                     := 'X';             -- wlast
			hps_0_h2f_lw_axi_master_wvalid                                      : in  std_logic                     := 'X';             -- wvalid
			hps_0_h2f_lw_axi_master_wready                                      : out std_logic;                                        -- wready
			hps_0_h2f_lw_axi_master_bid                                         : out std_logic_vector(11 downto 0);                    -- bid
			hps_0_h2f_lw_axi_master_bresp                                       : out std_logic_vector(1 downto 0);                     -- bresp
			hps_0_h2f_lw_axi_master_bvalid                                      : out std_logic;                                        -- bvalid
			hps_0_h2f_lw_axi_master_bready                                      : in  std_logic                     := 'X';             -- bready
			hps_0_h2f_lw_axi_master_arid                                        : in  std_logic_vector(11 downto 0) := (others => 'X'); -- arid
			hps_0_h2f_lw_axi_master_araddr                                      : in  std_logic_vector(20 downto 0) := (others => 'X'); -- araddr
			hps_0_h2f_lw_axi_master_arlen                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- arlen
			hps_0_h2f_lw_axi_master_arsize                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arsize
			hps_0_h2f_lw_axi_master_arburst                                     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- arburst
			hps_0_h2f_lw_axi_master_arlock                                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- arlock
			hps_0_h2f_lw_axi_master_arcache                                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- arcache
			hps_0_h2f_lw_axi_master_arprot                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arprot
			hps_0_h2f_lw_axi_master_arvalid                                     : in  std_logic                     := 'X';             -- arvalid
			hps_0_h2f_lw_axi_master_arready                                     : out std_logic;                                        -- arready
			hps_0_h2f_lw_axi_master_rid                                         : out std_logic_vector(11 downto 0);                    -- rid
			hps_0_h2f_lw_axi_master_rdata                                       : out std_logic_vector(31 downto 0);                    -- rdata
			hps_0_h2f_lw_axi_master_rresp                                       : out std_logic_vector(1 downto 0);                     -- rresp
			hps_0_h2f_lw_axi_master_rlast                                       : out std_logic;                                        -- rlast
			hps_0_h2f_lw_axi_master_rvalid                                      : out std_logic;                                        -- rvalid
			hps_0_h2f_lw_axi_master_rready                                      : in  std_logic                     := 'X';             -- rready
			clk_0_clk_clk                                                       : in  std_logic                     := 'X';             -- clk
			audio_0_reset_reset_bridge_in_reset_reset                           : in  std_logic                     := 'X';             -- reset
			hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			audio_0_avalon_audio_slave_address                                  : out std_logic_vector(1 downto 0);                     -- address
			audio_0_avalon_audio_slave_write                                    : out std_logic;                                        -- write
			audio_0_avalon_audio_slave_read                                     : out std_logic;                                        -- read
			audio_0_avalon_audio_slave_readdata                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			audio_0_avalon_audio_slave_writedata                                : out std_logic_vector(31 downto 0);                    -- writedata
			audio_0_avalon_audio_slave_chipselect                               : out std_logic;                                        -- chipselect
			audio_and_video_config_0_avalon_av_config_slave_address             : out std_logic_vector(1 downto 0);                     -- address
			audio_and_video_config_0_avalon_av_config_slave_write               : out std_logic;                                        -- write
			audio_and_video_config_0_avalon_av_config_slave_read                : out std_logic;                                        -- read
			audio_and_video_config_0_avalon_av_config_slave_readdata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			audio_and_video_config_0_avalon_av_config_slave_writedata           : out std_logic_vector(31 downto 0);                    -- writedata
			audio_and_video_config_0_avalon_av_config_slave_byteenable          : out std_logic_vector(3 downto 0);                     -- byteenable
			audio_and_video_config_0_avalon_av_config_slave_waitrequest         : in  std_logic                     := 'X';             -- waitrequest
			buttons_s1_address                                                  : out std_logic_vector(1 downto 0);                     -- address
			buttons_s1_write                                                    : out std_logic;                                        -- write
			buttons_s1_readdata                                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			buttons_s1_writedata                                                : out std_logic_vector(31 downto 0);                    -- writedata
			buttons_s1_chipselect                                               : out std_logic;                                        -- chipselect
			character_lcd_0_avalon_lcd_slave_address                            : out std_logic_vector(0 downto 0);                     -- address
			character_lcd_0_avalon_lcd_slave_write                              : out std_logic;                                        -- write
			character_lcd_0_avalon_lcd_slave_read                               : out std_logic;                                        -- read
			character_lcd_0_avalon_lcd_slave_readdata                           : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			character_lcd_0_avalon_lcd_slave_writedata                          : out std_logic_vector(7 downto 0);                     -- writedata
			character_lcd_0_avalon_lcd_slave_waitrequest                        : in  std_logic                     := 'X';             -- waitrequest
			character_lcd_0_avalon_lcd_slave_chipselect                         : out std_logic;                                        -- chipselect
			EnvelopeController_0_avalon_slave_write                             : out std_logic;                                        -- write
			EnvelopeController_0_avalon_slave_read                              : out std_logic;                                        -- read
			EnvelopeController_0_avalon_slave_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			EnvelopeController_0_avalon_slave_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			photodiode_0_avalon_slave_read                                      : out std_logic;                                        -- read
			photodiode_0_avalon_slave_readdata                                  : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			red_leds_s1_address                                                 : out std_logic_vector(1 downto 0);                     -- address
			red_leds_s1_write                                                   : out std_logic;                                        -- write
			red_leds_s1_readdata                                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			red_leds_s1_writedata                                               : out std_logic_vector(31 downto 0);                    -- writedata
			red_leds_s1_chipselect                                              : out std_logic;                                        -- chipselect
			switches_s1_address                                                 : out std_logic_vector(1 downto 0);                     -- address
			switches_s1_write                                                   : out std_logic;                                        -- write
			switches_s1_readdata                                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			switches_s1_writedata                                               : out std_logic_vector(31 downto 0);                    -- writedata
			switches_s1_chipselect                                              : out std_logic;                                        -- chipselect
			Synthesizer_0_avalon_slave_0_write                                  : out std_logic;                                        -- write
			Synthesizer_0_avalon_slave_0_read                                   : out std_logic;                                        -- read
			Synthesizer_0_avalon_slave_0_readdata                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Synthesizer_0_avalon_slave_0_writedata                              : out std_logic_vector(31 downto 0);                    -- writedata
			Synthesizer_1_avalon_slave_0_write                                  : out std_logic;                                        -- write
			Synthesizer_1_avalon_slave_0_read                                   : out std_logic;                                        -- read
			Synthesizer_1_avalon_slave_0_readdata                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Synthesizer_1_avalon_slave_0_writedata                              : out std_logic_vector(31 downto 0);                    -- writedata
			Synthesizer_2_avalon_slave_0_write                                  : out std_logic;                                        -- write
			Synthesizer_2_avalon_slave_0_read                                   : out std_logic;                                        -- read
			Synthesizer_2_avalon_slave_0_readdata                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Synthesizer_2_avalon_slave_0_writedata                              : out std_logic_vector(31 downto 0);                    -- writedata
			Synthesizer_3_avalon_slave_0_write                                  : out std_logic;                                        -- write
			Synthesizer_3_avalon_slave_0_read                                   : out std_logic;                                        -- read
			Synthesizer_3_avalon_slave_0_readdata                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Synthesizer_3_avalon_slave_0_writedata                              : out std_logic_vector(31 downto 0);                    -- writedata
			Synthesizer_4_avalon_slave_0_write                                  : out std_logic;                                        -- write
			Synthesizer_4_avalon_slave_0_read                                   : out std_logic;                                        -- read
			Synthesizer_4_avalon_slave_0_readdata                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Synthesizer_4_avalon_slave_0_writedata                              : out std_logic_vector(31 downto 0);                    -- writedata
			Synthesizer_5_avalon_slave_0_write                                  : out std_logic;                                        -- write
			Synthesizer_5_avalon_slave_0_read                                   : out std_logic;                                        -- read
			Synthesizer_5_avalon_slave_0_readdata                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Synthesizer_5_avalon_slave_0_writedata                              : out std_logic_vector(31 downto 0);                    -- writedata
			Synthesizer_6_avalon_slave_0_write                                  : out std_logic;                                        -- write
			Synthesizer_6_avalon_slave_0_read                                   : out std_logic;                                        -- read
			Synthesizer_6_avalon_slave_0_readdata                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Synthesizer_6_avalon_slave_0_writedata                              : out std_logic_vector(31 downto 0);                    -- writedata
			Synthesizer_7_avalon_slave_0_write                                  : out std_logic;                                        -- write
			Synthesizer_7_avalon_slave_0_read                                   : out std_logic;                                        -- read
			Synthesizer_7_avalon_slave_0_readdata                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Synthesizer_7_avalon_slave_0_writedata                              : out std_logic_vector(31 downto 0);                    -- writedata
			sysid_qsys_0_control_slave_address                                  : out std_logic_vector(0 downto 0);                     -- address
			sysid_qsys_0_control_slave_readdata                                 : in  std_logic_vector(31 downto 0) := (others => 'X')  -- readdata
		);
	end component soc_system_mm_interconnect_0;

	component soc_system_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component soc_system_irq_mapper;

	component soc_system_irq_mapper_001 is
		port (
			clk        : in  std_logic                     := 'X'; -- clk
			reset      : in  std_logic                     := 'X'; -- reset
			sender_irq : out std_logic_vector(31 downto 0)         -- irq
		);
	end component soc_system_irq_mapper_001;

	component soc_system_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component soc_system_rst_controller;

	component soc_system_rst_controller_002 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component soc_system_rst_controller_002;

	signal hps_0_h2f_lw_axi_master_awburst                                               : std_logic_vector(1 downto 0);  -- hps_0:h2f_lw_AWBURST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awburst
	signal hps_0_h2f_lw_axi_master_arlen                                                 : std_logic_vector(3 downto 0);  -- hps_0:h2f_lw_ARLEN -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arlen
	signal hps_0_h2f_lw_axi_master_wstrb                                                 : std_logic_vector(3 downto 0);  -- hps_0:h2f_lw_WSTRB -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wstrb
	signal hps_0_h2f_lw_axi_master_wready                                                : std_logic;                     -- mm_interconnect_0:hps_0_h2f_lw_axi_master_wready -> hps_0:h2f_lw_WREADY
	signal hps_0_h2f_lw_axi_master_rid                                                   : std_logic_vector(11 downto 0); -- mm_interconnect_0:hps_0_h2f_lw_axi_master_rid -> hps_0:h2f_lw_RID
	signal hps_0_h2f_lw_axi_master_rready                                                : std_logic;                     -- hps_0:h2f_lw_RREADY -> mm_interconnect_0:hps_0_h2f_lw_axi_master_rready
	signal hps_0_h2f_lw_axi_master_awlen                                                 : std_logic_vector(3 downto 0);  -- hps_0:h2f_lw_AWLEN -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awlen
	signal hps_0_h2f_lw_axi_master_wid                                                   : std_logic_vector(11 downto 0); -- hps_0:h2f_lw_WID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wid
	signal hps_0_h2f_lw_axi_master_arcache                                               : std_logic_vector(3 downto 0);  -- hps_0:h2f_lw_ARCACHE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arcache
	signal hps_0_h2f_lw_axi_master_wvalid                                                : std_logic;                     -- hps_0:h2f_lw_WVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wvalid
	signal hps_0_h2f_lw_axi_master_araddr                                                : std_logic_vector(20 downto 0); -- hps_0:h2f_lw_ARADDR -> mm_interconnect_0:hps_0_h2f_lw_axi_master_araddr
	signal hps_0_h2f_lw_axi_master_arprot                                                : std_logic_vector(2 downto 0);  -- hps_0:h2f_lw_ARPROT -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arprot
	signal hps_0_h2f_lw_axi_master_awprot                                                : std_logic_vector(2 downto 0);  -- hps_0:h2f_lw_AWPROT -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awprot
	signal hps_0_h2f_lw_axi_master_wdata                                                 : std_logic_vector(31 downto 0); -- hps_0:h2f_lw_WDATA -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wdata
	signal hps_0_h2f_lw_axi_master_arvalid                                               : std_logic;                     -- hps_0:h2f_lw_ARVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arvalid
	signal hps_0_h2f_lw_axi_master_awcache                                               : std_logic_vector(3 downto 0);  -- hps_0:h2f_lw_AWCACHE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awcache
	signal hps_0_h2f_lw_axi_master_arid                                                  : std_logic_vector(11 downto 0); -- hps_0:h2f_lw_ARID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arid
	signal hps_0_h2f_lw_axi_master_arlock                                                : std_logic_vector(1 downto 0);  -- hps_0:h2f_lw_ARLOCK -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arlock
	signal hps_0_h2f_lw_axi_master_awlock                                                : std_logic_vector(1 downto 0);  -- hps_0:h2f_lw_AWLOCK -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awlock
	signal hps_0_h2f_lw_axi_master_awaddr                                                : std_logic_vector(20 downto 0); -- hps_0:h2f_lw_AWADDR -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awaddr
	signal hps_0_h2f_lw_axi_master_bresp                                                 : std_logic_vector(1 downto 0);  -- mm_interconnect_0:hps_0_h2f_lw_axi_master_bresp -> hps_0:h2f_lw_BRESP
	signal hps_0_h2f_lw_axi_master_arready                                               : std_logic;                     -- mm_interconnect_0:hps_0_h2f_lw_axi_master_arready -> hps_0:h2f_lw_ARREADY
	signal hps_0_h2f_lw_axi_master_rdata                                                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:hps_0_h2f_lw_axi_master_rdata -> hps_0:h2f_lw_RDATA
	signal hps_0_h2f_lw_axi_master_awready                                               : std_logic;                     -- mm_interconnect_0:hps_0_h2f_lw_axi_master_awready -> hps_0:h2f_lw_AWREADY
	signal hps_0_h2f_lw_axi_master_arburst                                               : std_logic_vector(1 downto 0);  -- hps_0:h2f_lw_ARBURST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arburst
	signal hps_0_h2f_lw_axi_master_arsize                                                : std_logic_vector(2 downto 0);  -- hps_0:h2f_lw_ARSIZE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arsize
	signal hps_0_h2f_lw_axi_master_bready                                                : std_logic;                     -- hps_0:h2f_lw_BREADY -> mm_interconnect_0:hps_0_h2f_lw_axi_master_bready
	signal hps_0_h2f_lw_axi_master_rlast                                                 : std_logic;                     -- mm_interconnect_0:hps_0_h2f_lw_axi_master_rlast -> hps_0:h2f_lw_RLAST
	signal hps_0_h2f_lw_axi_master_wlast                                                 : std_logic;                     -- hps_0:h2f_lw_WLAST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wlast
	signal hps_0_h2f_lw_axi_master_rresp                                                 : std_logic_vector(1 downto 0);  -- mm_interconnect_0:hps_0_h2f_lw_axi_master_rresp -> hps_0:h2f_lw_RRESP
	signal hps_0_h2f_lw_axi_master_awid                                                  : std_logic_vector(11 downto 0); -- hps_0:h2f_lw_AWID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awid
	signal hps_0_h2f_lw_axi_master_bid                                                   : std_logic_vector(11 downto 0); -- mm_interconnect_0:hps_0_h2f_lw_axi_master_bid -> hps_0:h2f_lw_BID
	signal hps_0_h2f_lw_axi_master_bvalid                                                : std_logic;                     -- mm_interconnect_0:hps_0_h2f_lw_axi_master_bvalid -> hps_0:h2f_lw_BVALID
	signal hps_0_h2f_lw_axi_master_awsize                                                : std_logic_vector(2 downto 0);  -- hps_0:h2f_lw_AWSIZE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awsize
	signal hps_0_h2f_lw_axi_master_awvalid                                               : std_logic;                     -- hps_0:h2f_lw_AWVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awvalid
	signal hps_0_h2f_lw_axi_master_rvalid                                                : std_logic;                     -- mm_interconnect_0:hps_0_h2f_lw_axi_master_rvalid -> hps_0:h2f_lw_RVALID
	signal mm_interconnect_0_audio_0_avalon_audio_slave_chipselect                       : std_logic;                     -- mm_interconnect_0:audio_0_avalon_audio_slave_chipselect -> audio_0:chipselect
	signal mm_interconnect_0_audio_0_avalon_audio_slave_readdata                         : std_logic_vector(31 downto 0); -- audio_0:readdata -> mm_interconnect_0:audio_0_avalon_audio_slave_readdata
	signal mm_interconnect_0_audio_0_avalon_audio_slave_address                          : std_logic_vector(1 downto 0);  -- mm_interconnect_0:audio_0_avalon_audio_slave_address -> audio_0:address
	signal mm_interconnect_0_audio_0_avalon_audio_slave_read                             : std_logic;                     -- mm_interconnect_0:audio_0_avalon_audio_slave_read -> audio_0:read
	signal mm_interconnect_0_audio_0_avalon_audio_slave_write                            : std_logic;                     -- mm_interconnect_0:audio_0_avalon_audio_slave_write -> audio_0:write
	signal mm_interconnect_0_audio_0_avalon_audio_slave_writedata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:audio_0_avalon_audio_slave_writedata -> audio_0:writedata
	signal mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_readdata    : std_logic_vector(31 downto 0); -- audio_and_video_config_0:readdata -> mm_interconnect_0:audio_and_video_config_0_avalon_av_config_slave_readdata
	signal mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_waitrequest : std_logic;                     -- audio_and_video_config_0:waitrequest -> mm_interconnect_0:audio_and_video_config_0_avalon_av_config_slave_waitrequest
	signal mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_address     : std_logic_vector(1 downto 0);  -- mm_interconnect_0:audio_and_video_config_0_avalon_av_config_slave_address -> audio_and_video_config_0:address
	signal mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_read        : std_logic;                     -- mm_interconnect_0:audio_and_video_config_0_avalon_av_config_slave_read -> audio_and_video_config_0:read
	signal mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_byteenable  : std_logic_vector(3 downto 0);  -- mm_interconnect_0:audio_and_video_config_0_avalon_av_config_slave_byteenable -> audio_and_video_config_0:byteenable
	signal mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_write       : std_logic;                     -- mm_interconnect_0:audio_and_video_config_0_avalon_av_config_slave_write -> audio_and_video_config_0:write
	signal mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_writedata   : std_logic_vector(31 downto 0); -- mm_interconnect_0:audio_and_video_config_0_avalon_av_config_slave_writedata -> audio_and_video_config_0:writedata
	signal mm_interconnect_0_character_lcd_0_avalon_lcd_slave_chipselect                 : std_logic;                     -- mm_interconnect_0:character_lcd_0_avalon_lcd_slave_chipselect -> character_lcd_0:chipselect
	signal mm_interconnect_0_character_lcd_0_avalon_lcd_slave_readdata                   : std_logic_vector(7 downto 0);  -- character_lcd_0:readdata -> mm_interconnect_0:character_lcd_0_avalon_lcd_slave_readdata
	signal mm_interconnect_0_character_lcd_0_avalon_lcd_slave_waitrequest                : std_logic;                     -- character_lcd_0:waitrequest -> mm_interconnect_0:character_lcd_0_avalon_lcd_slave_waitrequest
	signal mm_interconnect_0_character_lcd_0_avalon_lcd_slave_address                    : std_logic_vector(0 downto 0);  -- mm_interconnect_0:character_lcd_0_avalon_lcd_slave_address -> character_lcd_0:address
	signal mm_interconnect_0_character_lcd_0_avalon_lcd_slave_read                       : std_logic;                     -- mm_interconnect_0:character_lcd_0_avalon_lcd_slave_read -> character_lcd_0:read
	signal mm_interconnect_0_character_lcd_0_avalon_lcd_slave_write                      : std_logic;                     -- mm_interconnect_0:character_lcd_0_avalon_lcd_slave_write -> character_lcd_0:write
	signal mm_interconnect_0_character_lcd_0_avalon_lcd_slave_writedata                  : std_logic_vector(7 downto 0);  -- mm_interconnect_0:character_lcd_0_avalon_lcd_slave_writedata -> character_lcd_0:writedata
	signal mm_interconnect_0_envelopecontroller_0_avalon_slave_readdata                  : std_logic_vector(31 downto 0); -- EnvelopeController_0:data_out -> mm_interconnect_0:EnvelopeController_0_avalon_slave_readdata
	signal mm_interconnect_0_envelopecontroller_0_avalon_slave_read                      : std_logic;                     -- mm_interconnect_0:EnvelopeController_0_avalon_slave_read -> EnvelopeController_0:read
	signal mm_interconnect_0_envelopecontroller_0_avalon_slave_write                     : std_logic;                     -- mm_interconnect_0:EnvelopeController_0_avalon_slave_write -> EnvelopeController_0:write
	signal mm_interconnect_0_envelopecontroller_0_avalon_slave_writedata                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:EnvelopeController_0_avalon_slave_writedata -> EnvelopeController_0:data_in
	signal mm_interconnect_0_photodiode_0_avalon_slave_readdata                          : std_logic_vector(7 downto 0);  -- photodiode_0:avalon_slave_readdata -> mm_interconnect_0:photodiode_0_avalon_slave_readdata
	signal mm_interconnect_0_photodiode_0_avalon_slave_read                              : std_logic;                     -- mm_interconnect_0:photodiode_0_avalon_slave_read -> mm_interconnect_0_photodiode_0_avalon_slave_read:in
	signal mm_interconnect_0_synthesizer_0_avalon_slave_0_readdata                       : std_logic_vector(31 downto 0); -- Synthesizer_0:data_out -> mm_interconnect_0:Synthesizer_0_avalon_slave_0_readdata
	signal mm_interconnect_0_synthesizer_0_avalon_slave_0_read                           : std_logic;                     -- mm_interconnect_0:Synthesizer_0_avalon_slave_0_read -> Synthesizer_0:read
	signal mm_interconnect_0_synthesizer_0_avalon_slave_0_write                          : std_logic;                     -- mm_interconnect_0:Synthesizer_0_avalon_slave_0_write -> Synthesizer_0:write
	signal mm_interconnect_0_synthesizer_0_avalon_slave_0_writedata                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:Synthesizer_0_avalon_slave_0_writedata -> Synthesizer_0:phase_reg
	signal mm_interconnect_0_synthesizer_1_avalon_slave_0_readdata                       : std_logic_vector(31 downto 0); -- Synthesizer_1:data_out -> mm_interconnect_0:Synthesizer_1_avalon_slave_0_readdata
	signal mm_interconnect_0_synthesizer_1_avalon_slave_0_read                           : std_logic;                     -- mm_interconnect_0:Synthesizer_1_avalon_slave_0_read -> Synthesizer_1:read
	signal mm_interconnect_0_synthesizer_1_avalon_slave_0_write                          : std_logic;                     -- mm_interconnect_0:Synthesizer_1_avalon_slave_0_write -> Synthesizer_1:write
	signal mm_interconnect_0_synthesizer_1_avalon_slave_0_writedata                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:Synthesizer_1_avalon_slave_0_writedata -> Synthesizer_1:phase_reg
	signal mm_interconnect_0_synthesizer_2_avalon_slave_0_readdata                       : std_logic_vector(31 downto 0); -- Synthesizer_2:data_out -> mm_interconnect_0:Synthesizer_2_avalon_slave_0_readdata
	signal mm_interconnect_0_synthesizer_2_avalon_slave_0_read                           : std_logic;                     -- mm_interconnect_0:Synthesizer_2_avalon_slave_0_read -> Synthesizer_2:read
	signal mm_interconnect_0_synthesizer_2_avalon_slave_0_write                          : std_logic;                     -- mm_interconnect_0:Synthesizer_2_avalon_slave_0_write -> Synthesizer_2:write
	signal mm_interconnect_0_synthesizer_2_avalon_slave_0_writedata                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:Synthesizer_2_avalon_slave_0_writedata -> Synthesizer_2:phase_reg
	signal mm_interconnect_0_synthesizer_3_avalon_slave_0_readdata                       : std_logic_vector(31 downto 0); -- Synthesizer_3:data_out -> mm_interconnect_0:Synthesizer_3_avalon_slave_0_readdata
	signal mm_interconnect_0_synthesizer_3_avalon_slave_0_read                           : std_logic;                     -- mm_interconnect_0:Synthesizer_3_avalon_slave_0_read -> Synthesizer_3:read
	signal mm_interconnect_0_synthesizer_3_avalon_slave_0_write                          : std_logic;                     -- mm_interconnect_0:Synthesizer_3_avalon_slave_0_write -> Synthesizer_3:write
	signal mm_interconnect_0_synthesizer_3_avalon_slave_0_writedata                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:Synthesizer_3_avalon_slave_0_writedata -> Synthesizer_3:phase_reg
	signal mm_interconnect_0_synthesizer_4_avalon_slave_0_readdata                       : std_logic_vector(31 downto 0); -- Synthesizer_4:data_out -> mm_interconnect_0:Synthesizer_4_avalon_slave_0_readdata
	signal mm_interconnect_0_synthesizer_4_avalon_slave_0_read                           : std_logic;                     -- mm_interconnect_0:Synthesizer_4_avalon_slave_0_read -> Synthesizer_4:read
	signal mm_interconnect_0_synthesizer_4_avalon_slave_0_write                          : std_logic;                     -- mm_interconnect_0:Synthesizer_4_avalon_slave_0_write -> Synthesizer_4:write
	signal mm_interconnect_0_synthesizer_4_avalon_slave_0_writedata                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:Synthesizer_4_avalon_slave_0_writedata -> Synthesizer_4:phase_reg
	signal mm_interconnect_0_synthesizer_5_avalon_slave_0_readdata                       : std_logic_vector(31 downto 0); -- Synthesizer_5:data_out -> mm_interconnect_0:Synthesizer_5_avalon_slave_0_readdata
	signal mm_interconnect_0_synthesizer_5_avalon_slave_0_read                           : std_logic;                     -- mm_interconnect_0:Synthesizer_5_avalon_slave_0_read -> Synthesizer_5:read
	signal mm_interconnect_0_synthesizer_5_avalon_slave_0_write                          : std_logic;                     -- mm_interconnect_0:Synthesizer_5_avalon_slave_0_write -> Synthesizer_5:write
	signal mm_interconnect_0_synthesizer_5_avalon_slave_0_writedata                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:Synthesizer_5_avalon_slave_0_writedata -> Synthesizer_5:phase_reg
	signal mm_interconnect_0_synthesizer_6_avalon_slave_0_readdata                       : std_logic_vector(31 downto 0); -- Synthesizer_6:data_out -> mm_interconnect_0:Synthesizer_6_avalon_slave_0_readdata
	signal mm_interconnect_0_synthesizer_6_avalon_slave_0_read                           : std_logic;                     -- mm_interconnect_0:Synthesizer_6_avalon_slave_0_read -> Synthesizer_6:read
	signal mm_interconnect_0_synthesizer_6_avalon_slave_0_write                          : std_logic;                     -- mm_interconnect_0:Synthesizer_6_avalon_slave_0_write -> Synthesizer_6:write
	signal mm_interconnect_0_synthesizer_6_avalon_slave_0_writedata                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:Synthesizer_6_avalon_slave_0_writedata -> Synthesizer_6:phase_reg
	signal mm_interconnect_0_synthesizer_7_avalon_slave_0_readdata                       : std_logic_vector(31 downto 0); -- Synthesizer_7:data_out -> mm_interconnect_0:Synthesizer_7_avalon_slave_0_readdata
	signal mm_interconnect_0_synthesizer_7_avalon_slave_0_read                           : std_logic;                     -- mm_interconnect_0:Synthesizer_7_avalon_slave_0_read -> Synthesizer_7:read
	signal mm_interconnect_0_synthesizer_7_avalon_slave_0_write                          : std_logic;                     -- mm_interconnect_0:Synthesizer_7_avalon_slave_0_write -> Synthesizer_7:write
	signal mm_interconnect_0_synthesizer_7_avalon_slave_0_writedata                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:Synthesizer_7_avalon_slave_0_writedata -> Synthesizer_7:phase_reg
	signal mm_interconnect_0_sysid_qsys_0_control_slave_readdata                         : std_logic_vector(31 downto 0); -- sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	signal mm_interconnect_0_sysid_qsys_0_control_slave_address                          : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	signal mm_interconnect_0_switches_s1_chipselect                                      : std_logic;                     -- mm_interconnect_0:switches_s1_chipselect -> switches:chipselect
	signal mm_interconnect_0_switches_s1_readdata                                        : std_logic_vector(31 downto 0); -- switches:readdata -> mm_interconnect_0:switches_s1_readdata
	signal mm_interconnect_0_switches_s1_address                                         : std_logic_vector(1 downto 0);  -- mm_interconnect_0:switches_s1_address -> switches:address
	signal mm_interconnect_0_switches_s1_write                                           : std_logic;                     -- mm_interconnect_0:switches_s1_write -> mm_interconnect_0_switches_s1_write:in
	signal mm_interconnect_0_switches_s1_writedata                                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:switches_s1_writedata -> switches:writedata
	signal mm_interconnect_0_buttons_s1_chipselect                                       : std_logic;                     -- mm_interconnect_0:buttons_s1_chipselect -> buttons:chipselect
	signal mm_interconnect_0_buttons_s1_readdata                                         : std_logic_vector(31 downto 0); -- buttons:readdata -> mm_interconnect_0:buttons_s1_readdata
	signal mm_interconnect_0_buttons_s1_address                                          : std_logic_vector(1 downto 0);  -- mm_interconnect_0:buttons_s1_address -> buttons:address
	signal mm_interconnect_0_buttons_s1_write                                            : std_logic;                     -- mm_interconnect_0:buttons_s1_write -> mm_interconnect_0_buttons_s1_write:in
	signal mm_interconnect_0_buttons_s1_writedata                                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:buttons_s1_writedata -> buttons:writedata
	signal mm_interconnect_0_red_leds_s1_chipselect                                      : std_logic;                     -- mm_interconnect_0:red_leds_s1_chipselect -> red_leds:chipselect
	signal mm_interconnect_0_red_leds_s1_readdata                                        : std_logic_vector(31 downto 0); -- red_leds:readdata -> mm_interconnect_0:red_leds_s1_readdata
	signal mm_interconnect_0_red_leds_s1_address                                         : std_logic_vector(1 downto 0);  -- mm_interconnect_0:red_leds_s1_address -> red_leds:address
	signal mm_interconnect_0_red_leds_s1_write                                           : std_logic;                     -- mm_interconnect_0:red_leds_s1_write -> mm_interconnect_0_red_leds_s1_write:in
	signal mm_interconnect_0_red_leds_s1_writedata                                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:red_leds_s1_writedata -> red_leds:writedata
	signal irq_mapper_receiver0_irq                                                      : std_logic;                     -- audio_0:irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                                      : std_logic;                     -- switches:irq -> irq_mapper:receiver1_irq
	signal irq_mapper_receiver2_irq                                                      : std_logic;                     -- buttons:irq -> irq_mapper:receiver2_irq
	signal hps_0_f2h_irq0_irq                                                            : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> hps_0:f2h_irq_p0
	signal hps_0_f2h_irq1_irq                                                            : std_logic_vector(31 downto 0); -- irq_mapper_001:sender_irq -> hps_0:f2h_irq_p1
	signal rst_controller_reset_out_reset                                                : std_logic;                     -- rst_controller:reset_out -> [EnvelopeController_0:reset, Synthesizer_0:reset, Synthesizer_1:reset, Synthesizer_2:reset, Synthesizer_3:reset, Synthesizer_4:reset, Synthesizer_5:reset, Synthesizer_6:reset, Synthesizer_7:reset, audio_0:reset, audio_and_video_config_0:reset, character_lcd_0:reset, mm_interconnect_0:audio_0_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in]
	signal hps_0_h2f_reset_reset                                                         : std_logic;                     -- hps_0:h2f_rst_n -> hps_0_h2f_reset_reset:in
	signal rst_controller_001_reset_out_reset                                            : std_logic;                     -- rst_controller_001:reset_out -> pll_0:rst
	signal rst_controller_002_reset_out_reset                                            : std_logic;                     -- rst_controller_002:reset_out -> mm_interconnect_0:hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset
	signal reset_reset_n_ports_inv                                                       : std_logic;                     -- reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0]
	signal mm_interconnect_0_photodiode_0_avalon_slave_read_ports_inv                    : std_logic;                     -- mm_interconnect_0_photodiode_0_avalon_slave_read:inv -> photodiode_0:avalon_slave_read_n
	signal mm_interconnect_0_switches_s1_write_ports_inv                                 : std_logic;                     -- mm_interconnect_0_switches_s1_write:inv -> switches:write_n
	signal mm_interconnect_0_buttons_s1_write_ports_inv                                  : std_logic;                     -- mm_interconnect_0_buttons_s1_write:inv -> buttons:write_n
	signal mm_interconnect_0_red_leds_s1_write_ports_inv                                 : std_logic;                     -- mm_interconnect_0_red_leds_s1_write:inv -> red_leds:write_n
	signal rst_controller_reset_out_reset_ports_inv                                      : std_logic;                     -- rst_controller_reset_out_reset:inv -> [buttons:reset_n, photodiode_0:reset_n, red_leds:reset_n, switches:reset_n, sysid_qsys_0:reset_n]
	signal hps_0_h2f_reset_reset_ports_inv                                               : std_logic;                     -- hps_0_h2f_reset_reset:inv -> [rst_controller:reset_in1, rst_controller_001:reset_in1, rst_controller_002:reset_in0]

begin

	envelopecontroller_0 : component EnvelopeController
		port map (
			data_out => mm_interconnect_0_envelopecontroller_0_avalon_slave_readdata,  -- avalon_slave.readdata
			read     => mm_interconnect_0_envelopecontroller_0_avalon_slave_read,      --             .read
			write    => mm_interconnect_0_envelopecontroller_0_avalon_slave_write,     --             .write
			data_in  => mm_interconnect_0_envelopecontroller_0_avalon_slave_writedata, --             .writedata
			reset    => rst_controller_reset_out_reset,                                --        reset.reset
			clk      => clk_clk                                                        --        clock.clk
		);

	synthesizer_0 : component synthesizer
		port map (
			clk       => clk_clk,                                                  --          clock.clk
			reset     => rst_controller_reset_out_reset,                           --          reset.reset
			phase_reg => mm_interconnect_0_synthesizer_0_avalon_slave_0_writedata, -- avalon_slave_0.writedata
			data_out  => mm_interconnect_0_synthesizer_0_avalon_slave_0_readdata,  --               .readdata
			read      => mm_interconnect_0_synthesizer_0_avalon_slave_0_read,      --               .read
			write     => mm_interconnect_0_synthesizer_0_avalon_slave_0_write      --               .write
		);

	synthesizer_1 : component synthesizer
		port map (
			clk       => clk_clk,                                                  --          clock.clk
			reset     => rst_controller_reset_out_reset,                           --          reset.reset
			phase_reg => mm_interconnect_0_synthesizer_1_avalon_slave_0_writedata, -- avalon_slave_0.writedata
			data_out  => mm_interconnect_0_synthesizer_1_avalon_slave_0_readdata,  --               .readdata
			read      => mm_interconnect_0_synthesizer_1_avalon_slave_0_read,      --               .read
			write     => mm_interconnect_0_synthesizer_1_avalon_slave_0_write      --               .write
		);

	synthesizer_2 : component synthesizer
		port map (
			clk       => clk_clk,                                                  --          clock.clk
			reset     => rst_controller_reset_out_reset,                           --          reset.reset
			phase_reg => mm_interconnect_0_synthesizer_2_avalon_slave_0_writedata, -- avalon_slave_0.writedata
			data_out  => mm_interconnect_0_synthesizer_2_avalon_slave_0_readdata,  --               .readdata
			read      => mm_interconnect_0_synthesizer_2_avalon_slave_0_read,      --               .read
			write     => mm_interconnect_0_synthesizer_2_avalon_slave_0_write      --               .write
		);

	synthesizer_3 : component synthesizer
		port map (
			clk       => clk_clk,                                                  --          clock.clk
			reset     => rst_controller_reset_out_reset,                           --          reset.reset
			phase_reg => mm_interconnect_0_synthesizer_3_avalon_slave_0_writedata, -- avalon_slave_0.writedata
			data_out  => mm_interconnect_0_synthesizer_3_avalon_slave_0_readdata,  --               .readdata
			read      => mm_interconnect_0_synthesizer_3_avalon_slave_0_read,      --               .read
			write     => mm_interconnect_0_synthesizer_3_avalon_slave_0_write      --               .write
		);

	synthesizer_4 : component synthesizer
		port map (
			clk       => clk_clk,                                                  --          clock.clk
			reset     => rst_controller_reset_out_reset,                           --          reset.reset
			phase_reg => mm_interconnect_0_synthesizer_4_avalon_slave_0_writedata, -- avalon_slave_0.writedata
			data_out  => mm_interconnect_0_synthesizer_4_avalon_slave_0_readdata,  --               .readdata
			read      => mm_interconnect_0_synthesizer_4_avalon_slave_0_read,      --               .read
			write     => mm_interconnect_0_synthesizer_4_avalon_slave_0_write      --               .write
		);

	synthesizer_5 : component synthesizer
		port map (
			clk       => clk_clk,                                                  --          clock.clk
			reset     => rst_controller_reset_out_reset,                           --          reset.reset
			phase_reg => mm_interconnect_0_synthesizer_5_avalon_slave_0_writedata, -- avalon_slave_0.writedata
			data_out  => mm_interconnect_0_synthesizer_5_avalon_slave_0_readdata,  --               .readdata
			read      => mm_interconnect_0_synthesizer_5_avalon_slave_0_read,      --               .read
			write     => mm_interconnect_0_synthesizer_5_avalon_slave_0_write      --               .write
		);

	synthesizer_6 : component synthesizer
		port map (
			clk       => clk_clk,                                                  --          clock.clk
			reset     => rst_controller_reset_out_reset,                           --          reset.reset
			phase_reg => mm_interconnect_0_synthesizer_6_avalon_slave_0_writedata, -- avalon_slave_0.writedata
			data_out  => mm_interconnect_0_synthesizer_6_avalon_slave_0_readdata,  --               .readdata
			read      => mm_interconnect_0_synthesizer_6_avalon_slave_0_read,      --               .read
			write     => mm_interconnect_0_synthesizer_6_avalon_slave_0_write      --               .write
		);

	synthesizer_7 : component synthesizer
		port map (
			clk       => clk_clk,                                                  --          clock.clk
			reset     => rst_controller_reset_out_reset,                           --          reset.reset
			phase_reg => mm_interconnect_0_synthesizer_7_avalon_slave_0_writedata, -- avalon_slave_0.writedata
			data_out  => mm_interconnect_0_synthesizer_7_avalon_slave_0_readdata,  --               .readdata
			read      => mm_interconnect_0_synthesizer_7_avalon_slave_0_read,      --               .read
			write     => mm_interconnect_0_synthesizer_7_avalon_slave_0_write      --               .write
		);

	audio_0 : component soc_system_audio_0
		port map (
			clk         => clk_clk,                                                 --                clk.clk
			reset       => rst_controller_reset_out_reset,                          --              reset.reset
			address     => mm_interconnect_0_audio_0_avalon_audio_slave_address,    -- avalon_audio_slave.address
			chipselect  => mm_interconnect_0_audio_0_avalon_audio_slave_chipselect, --                   .chipselect
			read        => mm_interconnect_0_audio_0_avalon_audio_slave_read,       --                   .read
			write       => mm_interconnect_0_audio_0_avalon_audio_slave_write,      --                   .write
			writedata   => mm_interconnect_0_audio_0_avalon_audio_slave_writedata,  --                   .writedata
			readdata    => mm_interconnect_0_audio_0_avalon_audio_slave_readdata,   --                   .readdata
			irq         => irq_mapper_receiver0_irq,                                --          interrupt.irq
			AUD_ADCDAT  => audio_0_external_interface_ADCDAT,                       -- external_interface.export
			AUD_ADCLRCK => audio_0_external_interface_ADCLRCK,                      --                   .export
			AUD_BCLK    => audio_0_external_interface_BCLK,                         --                   .export
			AUD_DACDAT  => audio_0_external_interface_DACDAT,                       --                   .export
			AUD_DACLRCK => audio_0_external_interface_DACLRCK                       --                   .export
		);

	audio_and_video_config_0 : component soc_system_audio_and_video_config_0
		port map (
			clk         => clk_clk,                                                                       --                    clk.clk
			reset       => rst_controller_reset_out_reset,                                                --                  reset.reset
			address     => mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_address,     -- avalon_av_config_slave.address
			byteenable  => mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_byteenable,  --                       .byteenable
			read        => mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_read,        --                       .read
			write       => mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_write,       --                       .write
			writedata   => mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_writedata,   --                       .writedata
			readdata    => mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_readdata,    --                       .readdata
			waitrequest => mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_waitrequest, --                       .waitrequest
			I2C_SDAT    => audio_and_video_config_0_external_interface_SDAT,                              --     external_interface.export
			I2C_SCLK    => audio_and_video_config_0_external_interface_SCLK                               --                       .export
		);

	buttons : component soc_system_buttons
		port map (
			clk        => clk_clk,                                      --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     --               reset.reset_n
			address    => mm_interconnect_0_buttons_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_buttons_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_buttons_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_buttons_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_buttons_s1_readdata,        --                    .readdata
			in_port    => buttons_external_connection_export,           -- external_connection.export
			irq        => irq_mapper_receiver2_irq                      --                 irq.irq
		);

	character_lcd_0 : component soc_system_character_lcd_0
		port map (
			clk         => clk_clk,                                                        --                clk.clk
			reset       => rst_controller_reset_out_reset,                                 --              reset.reset
			address     => mm_interconnect_0_character_lcd_0_avalon_lcd_slave_address(0),  --   avalon_lcd_slave.address
			chipselect  => mm_interconnect_0_character_lcd_0_avalon_lcd_slave_chipselect,  --                   .chipselect
			read        => mm_interconnect_0_character_lcd_0_avalon_lcd_slave_read,        --                   .read
			write       => mm_interconnect_0_character_lcd_0_avalon_lcd_slave_write,       --                   .write
			writedata   => mm_interconnect_0_character_lcd_0_avalon_lcd_slave_writedata,   --                   .writedata
			readdata    => mm_interconnect_0_character_lcd_0_avalon_lcd_slave_readdata,    --                   .readdata
			waitrequest => mm_interconnect_0_character_lcd_0_avalon_lcd_slave_waitrequest, --                   .waitrequest
			LCD_DATA    => character_lcd_0_external_interface_DATA,                        -- external_interface.export
			LCD_ON      => character_lcd_0_external_interface_ON,                          --                   .export
			LCD_BLON    => character_lcd_0_external_interface_BLON,                        --                   .export
			LCD_EN      => character_lcd_0_external_interface_EN,                          --                   .export
			LCD_RS      => character_lcd_0_external_interface_RS,                          --                   .export
			LCD_RW      => character_lcd_0_external_interface_RW                           --                   .export
		);

	hps_0 : component soc_system_hps_0
		generic map (
			F2S_Width => 0,
			S2F_Width => 0
		)
		port map (
			mem_a                    => memory_mem_a,                    --            memory.mem_a
			mem_ba                   => memory_mem_ba,                   --                  .mem_ba
			mem_ck                   => memory_mem_ck,                   --                  .mem_ck
			mem_ck_n                 => memory_mem_ck_n,                 --                  .mem_ck_n
			mem_cke                  => memory_mem_cke,                  --                  .mem_cke
			mem_cs_n                 => memory_mem_cs_n,                 --                  .mem_cs_n
			mem_ras_n                => memory_mem_ras_n,                --                  .mem_ras_n
			mem_cas_n                => memory_mem_cas_n,                --                  .mem_cas_n
			mem_we_n                 => memory_mem_we_n,                 --                  .mem_we_n
			mem_reset_n              => memory_mem_reset_n,              --                  .mem_reset_n
			mem_dq                   => memory_mem_dq,                   --                  .mem_dq
			mem_dqs                  => memory_mem_dqs,                  --                  .mem_dqs
			mem_dqs_n                => memory_mem_dqs_n,                --                  .mem_dqs_n
			mem_odt                  => memory_mem_odt,                  --                  .mem_odt
			mem_dm                   => memory_mem_dm,                   --                  .mem_dm
			oct_rzqin                => memory_oct_rzqin,                --                  .oct_rzqin
			hps_io_emac1_inst_TX_CLK => hps_io_hps_io_emac1_inst_TX_CLK, --            hps_io.hps_io_emac1_inst_TX_CLK
			hps_io_emac1_inst_TXD0   => hps_io_hps_io_emac1_inst_TXD0,   --                  .hps_io_emac1_inst_TXD0
			hps_io_emac1_inst_TXD1   => hps_io_hps_io_emac1_inst_TXD1,   --                  .hps_io_emac1_inst_TXD1
			hps_io_emac1_inst_TXD2   => hps_io_hps_io_emac1_inst_TXD2,   --                  .hps_io_emac1_inst_TXD2
			hps_io_emac1_inst_TXD3   => hps_io_hps_io_emac1_inst_TXD3,   --                  .hps_io_emac1_inst_TXD3
			hps_io_emac1_inst_RXD0   => hps_io_hps_io_emac1_inst_RXD0,   --                  .hps_io_emac1_inst_RXD0
			hps_io_emac1_inst_MDIO   => hps_io_hps_io_emac1_inst_MDIO,   --                  .hps_io_emac1_inst_MDIO
			hps_io_emac1_inst_MDC    => hps_io_hps_io_emac1_inst_MDC,    --                  .hps_io_emac1_inst_MDC
			hps_io_emac1_inst_RX_CTL => hps_io_hps_io_emac1_inst_RX_CTL, --                  .hps_io_emac1_inst_RX_CTL
			hps_io_emac1_inst_TX_CTL => hps_io_hps_io_emac1_inst_TX_CTL, --                  .hps_io_emac1_inst_TX_CTL
			hps_io_emac1_inst_RX_CLK => hps_io_hps_io_emac1_inst_RX_CLK, --                  .hps_io_emac1_inst_RX_CLK
			hps_io_emac1_inst_RXD1   => hps_io_hps_io_emac1_inst_RXD1,   --                  .hps_io_emac1_inst_RXD1
			hps_io_emac1_inst_RXD2   => hps_io_hps_io_emac1_inst_RXD2,   --                  .hps_io_emac1_inst_RXD2
			hps_io_emac1_inst_RXD3   => hps_io_hps_io_emac1_inst_RXD3,   --                  .hps_io_emac1_inst_RXD3
			hps_io_sdio_inst_CMD     => hps_io_hps_io_sdio_inst_CMD,     --                  .hps_io_sdio_inst_CMD
			hps_io_sdio_inst_D0      => hps_io_hps_io_sdio_inst_D0,      --                  .hps_io_sdio_inst_D0
			hps_io_sdio_inst_D1      => hps_io_hps_io_sdio_inst_D1,      --                  .hps_io_sdio_inst_D1
			hps_io_sdio_inst_CLK     => hps_io_hps_io_sdio_inst_CLK,     --                  .hps_io_sdio_inst_CLK
			hps_io_sdio_inst_D2      => hps_io_hps_io_sdio_inst_D2,      --                  .hps_io_sdio_inst_D2
			hps_io_sdio_inst_D3      => hps_io_hps_io_sdio_inst_D3,      --                  .hps_io_sdio_inst_D3
			hps_io_usb1_inst_D0      => hps_io_hps_io_usb1_inst_D0,      --                  .hps_io_usb1_inst_D0
			hps_io_usb1_inst_D1      => hps_io_hps_io_usb1_inst_D1,      --                  .hps_io_usb1_inst_D1
			hps_io_usb1_inst_D2      => hps_io_hps_io_usb1_inst_D2,      --                  .hps_io_usb1_inst_D2
			hps_io_usb1_inst_D3      => hps_io_hps_io_usb1_inst_D3,      --                  .hps_io_usb1_inst_D3
			hps_io_usb1_inst_D4      => hps_io_hps_io_usb1_inst_D4,      --                  .hps_io_usb1_inst_D4
			hps_io_usb1_inst_D5      => hps_io_hps_io_usb1_inst_D5,      --                  .hps_io_usb1_inst_D5
			hps_io_usb1_inst_D6      => hps_io_hps_io_usb1_inst_D6,      --                  .hps_io_usb1_inst_D6
			hps_io_usb1_inst_D7      => hps_io_hps_io_usb1_inst_D7,      --                  .hps_io_usb1_inst_D7
			hps_io_usb1_inst_CLK     => hps_io_hps_io_usb1_inst_CLK,     --                  .hps_io_usb1_inst_CLK
			hps_io_usb1_inst_STP     => hps_io_hps_io_usb1_inst_STP,     --                  .hps_io_usb1_inst_STP
			hps_io_usb1_inst_DIR     => hps_io_hps_io_usb1_inst_DIR,     --                  .hps_io_usb1_inst_DIR
			hps_io_usb1_inst_NXT     => hps_io_hps_io_usb1_inst_NXT,     --                  .hps_io_usb1_inst_NXT
			hps_io_spim1_inst_CLK    => hps_io_hps_io_spim1_inst_CLK,    --                  .hps_io_spim1_inst_CLK
			hps_io_spim1_inst_MOSI   => hps_io_hps_io_spim1_inst_MOSI,   --                  .hps_io_spim1_inst_MOSI
			hps_io_spim1_inst_MISO   => hps_io_hps_io_spim1_inst_MISO,   --                  .hps_io_spim1_inst_MISO
			hps_io_spim1_inst_SS0    => hps_io_hps_io_spim1_inst_SS0,    --                  .hps_io_spim1_inst_SS0
			hps_io_uart0_inst_RX     => hps_io_hps_io_uart0_inst_RX,     --                  .hps_io_uart0_inst_RX
			hps_io_uart0_inst_TX     => hps_io_hps_io_uart0_inst_TX,     --                  .hps_io_uart0_inst_TX
			hps_io_i2c0_inst_SDA     => hps_io_hps_io_i2c0_inst_SDA,     --                  .hps_io_i2c0_inst_SDA
			hps_io_i2c0_inst_SCL     => hps_io_hps_io_i2c0_inst_SCL,     --                  .hps_io_i2c0_inst_SCL
			hps_io_i2c1_inst_SDA     => hps_io_hps_io_i2c1_inst_SDA,     --                  .hps_io_i2c1_inst_SDA
			hps_io_i2c1_inst_SCL     => hps_io_hps_io_i2c1_inst_SCL,     --                  .hps_io_i2c1_inst_SCL
			hps_io_gpio_inst_GPIO09  => hps_io_hps_io_gpio_inst_GPIO09,  --                  .hps_io_gpio_inst_GPIO09
			hps_io_gpio_inst_GPIO35  => hps_io_hps_io_gpio_inst_GPIO35,  --                  .hps_io_gpio_inst_GPIO35
			hps_io_gpio_inst_GPIO40  => hps_io_hps_io_gpio_inst_GPIO40,  --                  .hps_io_gpio_inst_GPIO40
			hps_io_gpio_inst_GPIO48  => hps_io_hps_io_gpio_inst_GPIO48,  --                  .hps_io_gpio_inst_GPIO48
			hps_io_gpio_inst_GPIO53  => hps_io_hps_io_gpio_inst_GPIO53,  --                  .hps_io_gpio_inst_GPIO53
			hps_io_gpio_inst_GPIO54  => hps_io_hps_io_gpio_inst_GPIO54,  --                  .hps_io_gpio_inst_GPIO54
			hps_io_gpio_inst_GPIO61  => hps_io_hps_io_gpio_inst_GPIO61,  --                  .hps_io_gpio_inst_GPIO61
			h2f_rst_n                => hps_0_h2f_reset_reset,           --         h2f_reset.reset_n
			h2f_lw_axi_clk           => clk_clk,                         --  h2f_lw_axi_clock.clk
			h2f_lw_AWID              => hps_0_h2f_lw_axi_master_awid,    -- h2f_lw_axi_master.awid
			h2f_lw_AWADDR            => hps_0_h2f_lw_axi_master_awaddr,  --                  .awaddr
			h2f_lw_AWLEN             => hps_0_h2f_lw_axi_master_awlen,   --                  .awlen
			h2f_lw_AWSIZE            => hps_0_h2f_lw_axi_master_awsize,  --                  .awsize
			h2f_lw_AWBURST           => hps_0_h2f_lw_axi_master_awburst, --                  .awburst
			h2f_lw_AWLOCK            => hps_0_h2f_lw_axi_master_awlock,  --                  .awlock
			h2f_lw_AWCACHE           => hps_0_h2f_lw_axi_master_awcache, --                  .awcache
			h2f_lw_AWPROT            => hps_0_h2f_lw_axi_master_awprot,  --                  .awprot
			h2f_lw_AWVALID           => hps_0_h2f_lw_axi_master_awvalid, --                  .awvalid
			h2f_lw_AWREADY           => hps_0_h2f_lw_axi_master_awready, --                  .awready
			h2f_lw_WID               => hps_0_h2f_lw_axi_master_wid,     --                  .wid
			h2f_lw_WDATA             => hps_0_h2f_lw_axi_master_wdata,   --                  .wdata
			h2f_lw_WSTRB             => hps_0_h2f_lw_axi_master_wstrb,   --                  .wstrb
			h2f_lw_WLAST             => hps_0_h2f_lw_axi_master_wlast,   --                  .wlast
			h2f_lw_WVALID            => hps_0_h2f_lw_axi_master_wvalid,  --                  .wvalid
			h2f_lw_WREADY            => hps_0_h2f_lw_axi_master_wready,  --                  .wready
			h2f_lw_BID               => hps_0_h2f_lw_axi_master_bid,     --                  .bid
			h2f_lw_BRESP             => hps_0_h2f_lw_axi_master_bresp,   --                  .bresp
			h2f_lw_BVALID            => hps_0_h2f_lw_axi_master_bvalid,  --                  .bvalid
			h2f_lw_BREADY            => hps_0_h2f_lw_axi_master_bready,  --                  .bready
			h2f_lw_ARID              => hps_0_h2f_lw_axi_master_arid,    --                  .arid
			h2f_lw_ARADDR            => hps_0_h2f_lw_axi_master_araddr,  --                  .araddr
			h2f_lw_ARLEN             => hps_0_h2f_lw_axi_master_arlen,   --                  .arlen
			h2f_lw_ARSIZE            => hps_0_h2f_lw_axi_master_arsize,  --                  .arsize
			h2f_lw_ARBURST           => hps_0_h2f_lw_axi_master_arburst, --                  .arburst
			h2f_lw_ARLOCK            => hps_0_h2f_lw_axi_master_arlock,  --                  .arlock
			h2f_lw_ARCACHE           => hps_0_h2f_lw_axi_master_arcache, --                  .arcache
			h2f_lw_ARPROT            => hps_0_h2f_lw_axi_master_arprot,  --                  .arprot
			h2f_lw_ARVALID           => hps_0_h2f_lw_axi_master_arvalid, --                  .arvalid
			h2f_lw_ARREADY           => hps_0_h2f_lw_axi_master_arready, --                  .arready
			h2f_lw_RID               => hps_0_h2f_lw_axi_master_rid,     --                  .rid
			h2f_lw_RDATA             => hps_0_h2f_lw_axi_master_rdata,   --                  .rdata
			h2f_lw_RRESP             => hps_0_h2f_lw_axi_master_rresp,   --                  .rresp
			h2f_lw_RLAST             => hps_0_h2f_lw_axi_master_rlast,   --                  .rlast
			h2f_lw_RVALID            => hps_0_h2f_lw_axi_master_rvalid,  --                  .rvalid
			h2f_lw_RREADY            => hps_0_h2f_lw_axi_master_rready,  --                  .rready
			f2h_irq_p0               => hps_0_f2h_irq0_irq,              --          f2h_irq0.irq
			f2h_irq_p1               => hps_0_f2h_irq1_irq               --          f2h_irq1.irq
		);

	photodiode_0 : component photodiode
		port map (
			avalon_slave_readdata => mm_interconnect_0_photodiode_0_avalon_slave_readdata,       -- avalon_slave.readdata
			avalon_slave_read_n   => mm_interconnect_0_photodiode_0_avalon_slave_read_ports_inv, --             .read_n
			conduit_end_0         => photodiode_0_conduit_end_export0,                           --  conduit_end.export0
			conduit_end_1         => photodiode_0_conduit_end_export1,                           --             .export1
			conduit_end_2         => photodiode_0_conduit_end_export2,                           --             .export2
			conduit_end_3         => photodiode_0_conduit_end_export3,                           --             .export3
			conduit_end_4         => photodiode_0_conduit_end_export4,                           --             .export4
			conduit_end_5         => photodiode_0_conduit_end_export5,                           --             .export5
			conduit_end_6         => photodiode_0_conduit_end_export6,                           --             .export6
			conduit_end_7         => photodiode_0_conduit_end_export7,                           --             .export7
			clk                   => clk_clk,                                                    --        clock.clk
			reset_n               => rst_controller_reset_out_reset_ports_inv                    --        reset.reset_n
		);

	pll_0 : component soc_system_pll_0
		port map (
			refclk   => clk_clk,                            --  refclk.clk
			rst      => rst_controller_001_reset_out_reset, --   reset.reset
			outclk_0 => pll_0_outclk0_clk,                  -- outclk0.clk
			locked   => open                                -- (terminated)
		);

	red_leds : component soc_system_red_leds
		port map (
			clk        => clk_clk,                                       --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,      --               reset.reset_n
			address    => mm_interconnect_0_red_leds_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_red_leds_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_red_leds_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_red_leds_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_red_leds_s1_readdata,        --                    .readdata
			out_port   => red_leds_external_connection_export            -- external_connection.export
		);

	switches : component soc_system_switches
		port map (
			clk        => clk_clk,                                       --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,      --               reset.reset_n
			address    => mm_interconnect_0_switches_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_switches_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_switches_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_switches_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_switches_s1_readdata,        --                    .readdata
			in_port    => switches_external_connection_export,           -- external_connection.export
			irq        => irq_mapper_receiver1_irq                       --                 irq.irq
		);

	sysid_qsys_0 : component soc_system_sysid_qsys_0
		port map (
			clock    => clk_clk,                                                 --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,                --         reset.reset_n
			readdata => mm_interconnect_0_sysid_qsys_0_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_qsys_0_control_slave_address(0)  --              .address
		);

	mm_interconnect_0 : component soc_system_mm_interconnect_0
		port map (
			hps_0_h2f_lw_axi_master_awid                                        => hps_0_h2f_lw_axi_master_awid,                                                  --                                       hps_0_h2f_lw_axi_master.awid
			hps_0_h2f_lw_axi_master_awaddr                                      => hps_0_h2f_lw_axi_master_awaddr,                                                --                                                              .awaddr
			hps_0_h2f_lw_axi_master_awlen                                       => hps_0_h2f_lw_axi_master_awlen,                                                 --                                                              .awlen
			hps_0_h2f_lw_axi_master_awsize                                      => hps_0_h2f_lw_axi_master_awsize,                                                --                                                              .awsize
			hps_0_h2f_lw_axi_master_awburst                                     => hps_0_h2f_lw_axi_master_awburst,                                               --                                                              .awburst
			hps_0_h2f_lw_axi_master_awlock                                      => hps_0_h2f_lw_axi_master_awlock,                                                --                                                              .awlock
			hps_0_h2f_lw_axi_master_awcache                                     => hps_0_h2f_lw_axi_master_awcache,                                               --                                                              .awcache
			hps_0_h2f_lw_axi_master_awprot                                      => hps_0_h2f_lw_axi_master_awprot,                                                --                                                              .awprot
			hps_0_h2f_lw_axi_master_awvalid                                     => hps_0_h2f_lw_axi_master_awvalid,                                               --                                                              .awvalid
			hps_0_h2f_lw_axi_master_awready                                     => hps_0_h2f_lw_axi_master_awready,                                               --                                                              .awready
			hps_0_h2f_lw_axi_master_wid                                         => hps_0_h2f_lw_axi_master_wid,                                                   --                                                              .wid
			hps_0_h2f_lw_axi_master_wdata                                       => hps_0_h2f_lw_axi_master_wdata,                                                 --                                                              .wdata
			hps_0_h2f_lw_axi_master_wstrb                                       => hps_0_h2f_lw_axi_master_wstrb,                                                 --                                                              .wstrb
			hps_0_h2f_lw_axi_master_wlast                                       => hps_0_h2f_lw_axi_master_wlast,                                                 --                                                              .wlast
			hps_0_h2f_lw_axi_master_wvalid                                      => hps_0_h2f_lw_axi_master_wvalid,                                                --                                                              .wvalid
			hps_0_h2f_lw_axi_master_wready                                      => hps_0_h2f_lw_axi_master_wready,                                                --                                                              .wready
			hps_0_h2f_lw_axi_master_bid                                         => hps_0_h2f_lw_axi_master_bid,                                                   --                                                              .bid
			hps_0_h2f_lw_axi_master_bresp                                       => hps_0_h2f_lw_axi_master_bresp,                                                 --                                                              .bresp
			hps_0_h2f_lw_axi_master_bvalid                                      => hps_0_h2f_lw_axi_master_bvalid,                                                --                                                              .bvalid
			hps_0_h2f_lw_axi_master_bready                                      => hps_0_h2f_lw_axi_master_bready,                                                --                                                              .bready
			hps_0_h2f_lw_axi_master_arid                                        => hps_0_h2f_lw_axi_master_arid,                                                  --                                                              .arid
			hps_0_h2f_lw_axi_master_araddr                                      => hps_0_h2f_lw_axi_master_araddr,                                                --                                                              .araddr
			hps_0_h2f_lw_axi_master_arlen                                       => hps_0_h2f_lw_axi_master_arlen,                                                 --                                                              .arlen
			hps_0_h2f_lw_axi_master_arsize                                      => hps_0_h2f_lw_axi_master_arsize,                                                --                                                              .arsize
			hps_0_h2f_lw_axi_master_arburst                                     => hps_0_h2f_lw_axi_master_arburst,                                               --                                                              .arburst
			hps_0_h2f_lw_axi_master_arlock                                      => hps_0_h2f_lw_axi_master_arlock,                                                --                                                              .arlock
			hps_0_h2f_lw_axi_master_arcache                                     => hps_0_h2f_lw_axi_master_arcache,                                               --                                                              .arcache
			hps_0_h2f_lw_axi_master_arprot                                      => hps_0_h2f_lw_axi_master_arprot,                                                --                                                              .arprot
			hps_0_h2f_lw_axi_master_arvalid                                     => hps_0_h2f_lw_axi_master_arvalid,                                               --                                                              .arvalid
			hps_0_h2f_lw_axi_master_arready                                     => hps_0_h2f_lw_axi_master_arready,                                               --                                                              .arready
			hps_0_h2f_lw_axi_master_rid                                         => hps_0_h2f_lw_axi_master_rid,                                                   --                                                              .rid
			hps_0_h2f_lw_axi_master_rdata                                       => hps_0_h2f_lw_axi_master_rdata,                                                 --                                                              .rdata
			hps_0_h2f_lw_axi_master_rresp                                       => hps_0_h2f_lw_axi_master_rresp,                                                 --                                                              .rresp
			hps_0_h2f_lw_axi_master_rlast                                       => hps_0_h2f_lw_axi_master_rlast,                                                 --                                                              .rlast
			hps_0_h2f_lw_axi_master_rvalid                                      => hps_0_h2f_lw_axi_master_rvalid,                                                --                                                              .rvalid
			hps_0_h2f_lw_axi_master_rready                                      => hps_0_h2f_lw_axi_master_rready,                                                --                                                              .rready
			clk_0_clk_clk                                                       => clk_clk,                                                                       --                                                     clk_0_clk.clk
			audio_0_reset_reset_bridge_in_reset_reset                           => rst_controller_reset_out_reset,                                                --                           audio_0_reset_reset_bridge_in_reset.reset
			hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset => rst_controller_002_reset_out_reset,                                            -- hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
			audio_0_avalon_audio_slave_address                                  => mm_interconnect_0_audio_0_avalon_audio_slave_address,                          --                                    audio_0_avalon_audio_slave.address
			audio_0_avalon_audio_slave_write                                    => mm_interconnect_0_audio_0_avalon_audio_slave_write,                            --                                                              .write
			audio_0_avalon_audio_slave_read                                     => mm_interconnect_0_audio_0_avalon_audio_slave_read,                             --                                                              .read
			audio_0_avalon_audio_slave_readdata                                 => mm_interconnect_0_audio_0_avalon_audio_slave_readdata,                         --                                                              .readdata
			audio_0_avalon_audio_slave_writedata                                => mm_interconnect_0_audio_0_avalon_audio_slave_writedata,                        --                                                              .writedata
			audio_0_avalon_audio_slave_chipselect                               => mm_interconnect_0_audio_0_avalon_audio_slave_chipselect,                       --                                                              .chipselect
			audio_and_video_config_0_avalon_av_config_slave_address             => mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_address,     --               audio_and_video_config_0_avalon_av_config_slave.address
			audio_and_video_config_0_avalon_av_config_slave_write               => mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_write,       --                                                              .write
			audio_and_video_config_0_avalon_av_config_slave_read                => mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_read,        --                                                              .read
			audio_and_video_config_0_avalon_av_config_slave_readdata            => mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_readdata,    --                                                              .readdata
			audio_and_video_config_0_avalon_av_config_slave_writedata           => mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_writedata,   --                                                              .writedata
			audio_and_video_config_0_avalon_av_config_slave_byteenable          => mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_byteenable,  --                                                              .byteenable
			audio_and_video_config_0_avalon_av_config_slave_waitrequest         => mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_waitrequest, --                                                              .waitrequest
			buttons_s1_address                                                  => mm_interconnect_0_buttons_s1_address,                                          --                                                    buttons_s1.address
			buttons_s1_write                                                    => mm_interconnect_0_buttons_s1_write,                                            --                                                              .write
			buttons_s1_readdata                                                 => mm_interconnect_0_buttons_s1_readdata,                                         --                                                              .readdata
			buttons_s1_writedata                                                => mm_interconnect_0_buttons_s1_writedata,                                        --                                                              .writedata
			buttons_s1_chipselect                                               => mm_interconnect_0_buttons_s1_chipselect,                                       --                                                              .chipselect
			character_lcd_0_avalon_lcd_slave_address                            => mm_interconnect_0_character_lcd_0_avalon_lcd_slave_address,                    --                              character_lcd_0_avalon_lcd_slave.address
			character_lcd_0_avalon_lcd_slave_write                              => mm_interconnect_0_character_lcd_0_avalon_lcd_slave_write,                      --                                                              .write
			character_lcd_0_avalon_lcd_slave_read                               => mm_interconnect_0_character_lcd_0_avalon_lcd_slave_read,                       --                                                              .read
			character_lcd_0_avalon_lcd_slave_readdata                           => mm_interconnect_0_character_lcd_0_avalon_lcd_slave_readdata,                   --                                                              .readdata
			character_lcd_0_avalon_lcd_slave_writedata                          => mm_interconnect_0_character_lcd_0_avalon_lcd_slave_writedata,                  --                                                              .writedata
			character_lcd_0_avalon_lcd_slave_waitrequest                        => mm_interconnect_0_character_lcd_0_avalon_lcd_slave_waitrequest,                --                                                              .waitrequest
			character_lcd_0_avalon_lcd_slave_chipselect                         => mm_interconnect_0_character_lcd_0_avalon_lcd_slave_chipselect,                 --                                                              .chipselect
			EnvelopeController_0_avalon_slave_write                             => mm_interconnect_0_envelopecontroller_0_avalon_slave_write,                     --                             EnvelopeController_0_avalon_slave.write
			EnvelopeController_0_avalon_slave_read                              => mm_interconnect_0_envelopecontroller_0_avalon_slave_read,                      --                                                              .read
			EnvelopeController_0_avalon_slave_readdata                          => mm_interconnect_0_envelopecontroller_0_avalon_slave_readdata,                  --                                                              .readdata
			EnvelopeController_0_avalon_slave_writedata                         => mm_interconnect_0_envelopecontroller_0_avalon_slave_writedata,                 --                                                              .writedata
			photodiode_0_avalon_slave_read                                      => mm_interconnect_0_photodiode_0_avalon_slave_read,                              --                                     photodiode_0_avalon_slave.read
			photodiode_0_avalon_slave_readdata                                  => mm_interconnect_0_photodiode_0_avalon_slave_readdata,                          --                                                              .readdata
			red_leds_s1_address                                                 => mm_interconnect_0_red_leds_s1_address,                                         --                                                   red_leds_s1.address
			red_leds_s1_write                                                   => mm_interconnect_0_red_leds_s1_write,                                           --                                                              .write
			red_leds_s1_readdata                                                => mm_interconnect_0_red_leds_s1_readdata,                                        --                                                              .readdata
			red_leds_s1_writedata                                               => mm_interconnect_0_red_leds_s1_writedata,                                       --                                                              .writedata
			red_leds_s1_chipselect                                              => mm_interconnect_0_red_leds_s1_chipselect,                                      --                                                              .chipselect
			switches_s1_address                                                 => mm_interconnect_0_switches_s1_address,                                         --                                                   switches_s1.address
			switches_s1_write                                                   => mm_interconnect_0_switches_s1_write,                                           --                                                              .write
			switches_s1_readdata                                                => mm_interconnect_0_switches_s1_readdata,                                        --                                                              .readdata
			switches_s1_writedata                                               => mm_interconnect_0_switches_s1_writedata,                                       --                                                              .writedata
			switches_s1_chipselect                                              => mm_interconnect_0_switches_s1_chipselect,                                      --                                                              .chipselect
			Synthesizer_0_avalon_slave_0_write                                  => mm_interconnect_0_synthesizer_0_avalon_slave_0_write,                          --                                  Synthesizer_0_avalon_slave_0.write
			Synthesizer_0_avalon_slave_0_read                                   => mm_interconnect_0_synthesizer_0_avalon_slave_0_read,                           --                                                              .read
			Synthesizer_0_avalon_slave_0_readdata                               => mm_interconnect_0_synthesizer_0_avalon_slave_0_readdata,                       --                                                              .readdata
			Synthesizer_0_avalon_slave_0_writedata                              => mm_interconnect_0_synthesizer_0_avalon_slave_0_writedata,                      --                                                              .writedata
			Synthesizer_1_avalon_slave_0_write                                  => mm_interconnect_0_synthesizer_1_avalon_slave_0_write,                          --                                  Synthesizer_1_avalon_slave_0.write
			Synthesizer_1_avalon_slave_0_read                                   => mm_interconnect_0_synthesizer_1_avalon_slave_0_read,                           --                                                              .read
			Synthesizer_1_avalon_slave_0_readdata                               => mm_interconnect_0_synthesizer_1_avalon_slave_0_readdata,                       --                                                              .readdata
			Synthesizer_1_avalon_slave_0_writedata                              => mm_interconnect_0_synthesizer_1_avalon_slave_0_writedata,                      --                                                              .writedata
			Synthesizer_2_avalon_slave_0_write                                  => mm_interconnect_0_synthesizer_2_avalon_slave_0_write,                          --                                  Synthesizer_2_avalon_slave_0.write
			Synthesizer_2_avalon_slave_0_read                                   => mm_interconnect_0_synthesizer_2_avalon_slave_0_read,                           --                                                              .read
			Synthesizer_2_avalon_slave_0_readdata                               => mm_interconnect_0_synthesizer_2_avalon_slave_0_readdata,                       --                                                              .readdata
			Synthesizer_2_avalon_slave_0_writedata                              => mm_interconnect_0_synthesizer_2_avalon_slave_0_writedata,                      --                                                              .writedata
			Synthesizer_3_avalon_slave_0_write                                  => mm_interconnect_0_synthesizer_3_avalon_slave_0_write,                          --                                  Synthesizer_3_avalon_slave_0.write
			Synthesizer_3_avalon_slave_0_read                                   => mm_interconnect_0_synthesizer_3_avalon_slave_0_read,                           --                                                              .read
			Synthesizer_3_avalon_slave_0_readdata                               => mm_interconnect_0_synthesizer_3_avalon_slave_0_readdata,                       --                                                              .readdata
			Synthesizer_3_avalon_slave_0_writedata                              => mm_interconnect_0_synthesizer_3_avalon_slave_0_writedata,                      --                                                              .writedata
			Synthesizer_4_avalon_slave_0_write                                  => mm_interconnect_0_synthesizer_4_avalon_slave_0_write,                          --                                  Synthesizer_4_avalon_slave_0.write
			Synthesizer_4_avalon_slave_0_read                                   => mm_interconnect_0_synthesizer_4_avalon_slave_0_read,                           --                                                              .read
			Synthesizer_4_avalon_slave_0_readdata                               => mm_interconnect_0_synthesizer_4_avalon_slave_0_readdata,                       --                                                              .readdata
			Synthesizer_4_avalon_slave_0_writedata                              => mm_interconnect_0_synthesizer_4_avalon_slave_0_writedata,                      --                                                              .writedata
			Synthesizer_5_avalon_slave_0_write                                  => mm_interconnect_0_synthesizer_5_avalon_slave_0_write,                          --                                  Synthesizer_5_avalon_slave_0.write
			Synthesizer_5_avalon_slave_0_read                                   => mm_interconnect_0_synthesizer_5_avalon_slave_0_read,                           --                                                              .read
			Synthesizer_5_avalon_slave_0_readdata                               => mm_interconnect_0_synthesizer_5_avalon_slave_0_readdata,                       --                                                              .readdata
			Synthesizer_5_avalon_slave_0_writedata                              => mm_interconnect_0_synthesizer_5_avalon_slave_0_writedata,                      --                                                              .writedata
			Synthesizer_6_avalon_slave_0_write                                  => mm_interconnect_0_synthesizer_6_avalon_slave_0_write,                          --                                  Synthesizer_6_avalon_slave_0.write
			Synthesizer_6_avalon_slave_0_read                                   => mm_interconnect_0_synthesizer_6_avalon_slave_0_read,                           --                                                              .read
			Synthesizer_6_avalon_slave_0_readdata                               => mm_interconnect_0_synthesizer_6_avalon_slave_0_readdata,                       --                                                              .readdata
			Synthesizer_6_avalon_slave_0_writedata                              => mm_interconnect_0_synthesizer_6_avalon_slave_0_writedata,                      --                                                              .writedata
			Synthesizer_7_avalon_slave_0_write                                  => mm_interconnect_0_synthesizer_7_avalon_slave_0_write,                          --                                  Synthesizer_7_avalon_slave_0.write
			Synthesizer_7_avalon_slave_0_read                                   => mm_interconnect_0_synthesizer_7_avalon_slave_0_read,                           --                                                              .read
			Synthesizer_7_avalon_slave_0_readdata                               => mm_interconnect_0_synthesizer_7_avalon_slave_0_readdata,                       --                                                              .readdata
			Synthesizer_7_avalon_slave_0_writedata                              => mm_interconnect_0_synthesizer_7_avalon_slave_0_writedata,                      --                                                              .writedata
			sysid_qsys_0_control_slave_address                                  => mm_interconnect_0_sysid_qsys_0_control_slave_address,                          --                                    sysid_qsys_0_control_slave.address
			sysid_qsys_0_control_slave_readdata                                 => mm_interconnect_0_sysid_qsys_0_control_slave_readdata                          --                                                              .readdata
		);

	irq_mapper : component soc_system_irq_mapper
		port map (
			clk           => open,                     --       clk.clk
			reset         => open,                     -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq, -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq, -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq, -- receiver2.irq
			sender_irq    => hps_0_f2h_irq0_irq        --    sender.irq
		);

	irq_mapper_001 : component soc_system_irq_mapper_001
		port map (
			clk        => open,               --       clk.clk
			reset      => open,               -- clk_reset.reset
			sender_irq => hps_0_f2h_irq1_irq  --    sender.irq
		);

	rst_controller : component soc_system_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,         -- reset_in0.reset
			reset_in1      => hps_0_h2f_reset_reset_ports_inv, -- reset_in1.reset
			clk            => clk_clk,                         --       clk.clk
			reset_out      => rst_controller_reset_out_reset,  -- reset_out.reset
			reset_req      => open,                            -- (terminated)
			reset_req_in0  => '0',                             -- (terminated)
			reset_req_in1  => '0',                             -- (terminated)
			reset_in2      => '0',                             -- (terminated)
			reset_req_in2  => '0',                             -- (terminated)
			reset_in3      => '0',                             -- (terminated)
			reset_req_in3  => '0',                             -- (terminated)
			reset_in4      => '0',                             -- (terminated)
			reset_req_in4  => '0',                             -- (terminated)
			reset_in5      => '0',                             -- (terminated)
			reset_req_in5  => '0',                             -- (terminated)
			reset_in6      => '0',                             -- (terminated)
			reset_req_in6  => '0',                             -- (terminated)
			reset_in7      => '0',                             -- (terminated)
			reset_req_in7  => '0',                             -- (terminated)
			reset_in8      => '0',                             -- (terminated)
			reset_req_in8  => '0',                             -- (terminated)
			reset_in9      => '0',                             -- (terminated)
			reset_req_in9  => '0',                             -- (terminated)
			reset_in10     => '0',                             -- (terminated)
			reset_req_in10 => '0',                             -- (terminated)
			reset_in11     => '0',                             -- (terminated)
			reset_req_in11 => '0',                             -- (terminated)
			reset_in12     => '0',                             -- (terminated)
			reset_req_in12 => '0',                             -- (terminated)
			reset_in13     => '0',                             -- (terminated)
			reset_req_in13 => '0',                             -- (terminated)
			reset_in14     => '0',                             -- (terminated)
			reset_req_in14 => '0',                             -- (terminated)
			reset_in15     => '0',                             -- (terminated)
			reset_req_in15 => '0'                              -- (terminated)
		);

	rst_controller_001 : component soc_system_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "none",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			reset_in1      => hps_0_h2f_reset_reset_ports_inv,    -- reset_in1.reset
			clk            => open,                               --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_002 : component soc_system_rst_controller_002
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => hps_0_h2f_reset_reset_ports_inv,    -- reset_in0.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_002_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_photodiode_0_avalon_slave_read_ports_inv <= not mm_interconnect_0_photodiode_0_avalon_slave_read;

	mm_interconnect_0_switches_s1_write_ports_inv <= not mm_interconnect_0_switches_s1_write;

	mm_interconnect_0_buttons_s1_write_ports_inv <= not mm_interconnect_0_buttons_s1_write;

	mm_interconnect_0_red_leds_s1_write_ports_inv <= not mm_interconnect_0_red_leds_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	hps_0_h2f_reset_reset_ports_inv <= not hps_0_h2f_reset_reset;

end architecture rtl; -- of soc_system
