 --------------------------------------------------------------------------------------------------------------------------
-- Original Authors : Simon Doherty, Eric Lunty, Kyle Brooks, Peter Roland						--
-- Date created: N/A 													--
--															--
-- Additional Authors : Randi Derbyshire, Adam Narten, Oliver Rarog, Celeste Chiasson					--
-- Date edited: March 26, 2018											--
--															--
-- This program takes a value from the synthesizer.vhd file and runs it through the 12-bit ROM to find the 	 	--
-- respective sine wave value. 												--
--------------------------------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use IEEE.STD_LOGIC_SIGNED.all;
use ieee.numeric_std.all;               -- Needed for shifts

entity HarpsichordSin_lut is

port (
	clk      : in  std_logic;
	en       : in  std_logic;
	
	--Address input
	address_reg : in std_logic_vector(11 downto 0); 
	
	--Sine value output
	sin_out  : out std_logic_vector(31 downto 0)
	);
end entity;


architecture rtl of HarpsichordSin_lut is


type rom_type is array (0 to 4095) of std_logic_vector (11 downto 0);

constant SIN_ROM : rom_type :=

(
X"86D", X"86F", X"871", X"873", X"876", X"878", X"87A", X"87C", 
X"87E", X"880", X"882", X"884", X"887", X"889", X"88B", X"88D", 
X"88F", X"891", X"894", X"896", X"898", X"89A", X"89C", X"89E", 
X"8A0", X"8A3", X"8A5", X"8A7", X"8A9", X"8AB", X"8AD", X"8B0", 
X"8B2", X"8B4", X"8B6", X"8B8", X"8BA", X"8BC", X"8BE", X"8C1", 
X"8C3", X"8C5", X"8C7", X"8C9", X"8CB", X"8CD", X"8D0", X"8D2", 
X"8D4", X"8D6", X"8D8", X"8DA", X"8DD", X"8DF", X"8E1", X"8E3", 
X"8E5", X"8E7", X"8E9", X"8EB", X"8EE", X"8F0", X"8F2", X"8F4", 
X"8F6", X"8F8", X"8FB", X"8FD", X"8FF", X"901", X"903", X"905", 
X"907", X"90A", X"90C", X"90E", X"910", X"912", X"914", X"916", 
X"918", X"91B", X"91D", X"91F", X"921", X"923", X"925", X"928", 
X"92A", X"92C", X"92E", X"930", X"932", X"934", X"937", X"939", 
X"93B", X"93D", X"93F", X"941", X"943", X"945", X"948", X"94A", 
X"94C", X"94E", X"950", X"952", X"955", X"957", X"959", X"95B", 
X"95D", X"95F", X"961", X"964", X"966", X"968", X"96A", X"96C", 
X"96E", X"970", X"973", X"975", X"977", X"979", X"97B", X"97D", 
X"97F", X"982", X"984", X"986", X"988", X"98A", X"98C", X"98E", 
X"991", X"993", X"995", X"997", X"999", X"99B", X"99D", X"9A0", 
X"9A2", X"9A4", X"9A6", X"9A8", X"9AA", X"9AC", X"9AF", X"9B1", 
X"9B3", X"9B5", X"9B7", X"9B9", X"9BC", X"9BE", X"9C0", X"9C2", 
X"9C4", X"9C6", X"9C8", X"9CA", X"9CD", X"9CF", X"9D1", X"9D3", 
X"9D5", X"9D7", X"9D9", X"9DC", X"9DE", X"9E0", X"9E2", X"9E4", 
X"9E6", X"9E9", X"9EB", X"9ED", X"9EF", X"9F1", X"9F3", X"9F5", 
X"9F7", X"9FA", X"9FC", X"9FE", X"A00", X"A02", X"A04", X"A06", 
X"A09", X"A0B", X"A0D", X"A0F", X"A11", X"A13", X"A16", X"A18", 
X"A1A", X"A1C", X"A1E", X"A20", X"A22", X"A24", X"A27", X"A29", 
X"A2B", X"A2D", X"A2F", X"A31", X"A34", X"A36", X"A38", X"A3A", 
X"A3C", X"A3E", X"A40", X"A43", X"A45", X"A47", X"A49", X"A4B", 
X"A4D", X"A4F", X"A51", X"A54", X"A56", X"A58", X"A5A", X"A5C", 
X"A5E", X"A61", X"A63", X"A65", X"A67", X"A69", X"A6B", X"A6D", 
X"A70", X"A72", X"A74", X"A76", X"A78", X"A7A", X"A7C", X"A7E", 
X"A81", X"A83", X"A85", X"A87", X"A89", X"A8B", X"A8E", X"A90", 
X"A92", X"A94", X"A96", X"A98", X"A9A", X"A9D", X"A9F", X"AA1", 
X"AA3", X"AA5", X"AA7", X"AA9", X"AAB", X"AAE", X"AB0", X"AB2", 
X"AB4", X"AB6", X"AB8", X"ABB", X"ABD", X"ABF", X"AC1", X"AC3", 
X"AC5", X"AC7", X"ACA", X"ACC", X"ACE", X"AD0", X"AD2", X"AD4", 
X"AD6", X"AD9", X"ADB", X"ADD", X"ADF", X"AE1", X"AE3", X"AE5", 
X"AE8", X"AEA", X"AEC", X"AEE", X"AF0", X"AF2", X"AF5", X"AF7", 
X"AF9", X"AFB", X"AFD", X"AFF", X"B01", X"B03", X"B06", X"B08", 
X"B0A", X"B0C", X"B0E", X"B10", X"B12", X"B15", X"B17", X"B19", 
X"B1B", X"B1D", X"B1F", X"B22", X"B24", X"B26", X"B28", X"B2A", 
X"B2C", X"B2E", X"B30", X"B33", X"B35", X"B37", X"B39", X"B3B", 
X"B3D", X"B3F", X"B42", X"B44", X"B46", X"B48", X"B4A", X"B4C", 
X"B4F", X"B51", X"B53", X"B55", X"B57", X"B59", X"B5B", X"B5E", 
X"B60", X"B62", X"B64", X"B66", X"B68", X"B6A", X"B6C", X"B6F", 
X"B71", X"B73", X"B75", X"B77", X"B79", X"B7C", X"B7E", X"B80", 
X"B82", X"B84", X"B86", X"B88", X"B8B", X"B8D", X"B8F", X"B91", 
X"B93", X"B95", X"B97", X"B9A", X"B9C", X"B9E", X"BA0", X"BA2", 
X"BA4", X"BA6", X"BA9", X"BAB", X"BAD", X"BAF", X"BB1", X"BB3", 
X"BB6", X"BB8", X"BBA", X"BBC", X"BBE", X"BC0", X"BC2", X"BC4", 
X"BC7", X"BC9", X"BCB", X"BCD", X"BCF", X"BD1", X"BD3", X"BD6", 
X"BD8", X"BDA", X"BDC", X"BDE", X"BE0", X"BE3", X"BE5", X"BE7", 
X"BE9", X"BEB", X"BED", X"BEF", X"BF1", X"BF4", X"BF6", X"BF8", 
X"BFA", X"BFC", X"BFE", X"C00", X"C03", X"C05", X"C07", X"C09", 
X"C0B", X"C0D", X"C10", X"C12", X"C14", X"C16", X"C18", X"C1A", 
X"C1C", X"C1E", X"C21", X"C23", X"C25", X"C27", X"C29", X"C2B", 
X"C2D", X"C30", X"C32", X"C34", X"C36", X"C38", X"C3A", X"C3D", 
X"C3F", X"C41", X"C43", X"C45", X"C47", X"C49", X"C4B", X"C4E", 
X"C50", X"C52", X"C54", X"C56", X"C58", X"C5B", X"C5D", X"C5F", 
X"C61", X"C63", X"C65", X"C67", X"C6A", X"C6C", X"C6E", X"C70", 
X"C72", X"C74", X"C76", X"C78", X"C7B", X"C7D", X"C7F", X"C81", 
X"C83", X"C85", X"C88", X"C8A", X"C8C", X"C8E", X"C90", X"C92", 
X"C94", X"C97", X"C99", X"C9B", X"C9D", X"C9F", X"CA1", X"CA3", 
X"CA5", X"CA8", X"CAA", X"CAC", X"CAE", X"CB0", X"CB2", X"CB5", 
X"CB7", X"CB9", X"CBB", X"CBD", X"CBF", X"CC1", X"CC4", X"CC6", 
X"CC8", X"CCA", X"CCC", X"CCE", X"CD0", X"CD2", X"CD5", X"CD7", 
X"CD9", X"CDB", X"CDD", X"CDF", X"CE2", X"CE4", X"CE6", X"CE8", 
X"CEA", X"CEC", X"CEE", X"CF1", X"CF3", X"CF5", X"CF7", X"CF9", 
X"CFB", X"CFD", X"D00", X"D02", X"D04", X"D06", X"D08", X"D0A", 
X"D0C", X"D0F", X"D11", X"D13", X"D15", X"D17", X"D19", X"D1C", 
X"D1E", X"D20", X"D22", X"D24", X"D26", X"D28", X"D2A", X"D2D", 
X"D2F", X"D31", X"D33", X"D35", X"D37", X"D39", X"D3C", X"D3E", 
X"D40", X"D42", X"D44", X"D46", X"D49", X"D4B", X"D4D", X"D4F", 
X"D51", X"D53", X"D41", X"D43", X"D45", X"D47", X"D49", X"D4C", 
X"D4E", X"D50", X"D52", X"D54", X"D56", X"D59", X"D5B", X"D5D", 
X"D5F", X"D61", X"D63", X"D65", X"D67", X"D6A", X"D6C", X"D6E", 
X"D70", X"D72", X"D74", X"D76", X"D79", X"D7B", X"D7D", X"D7F", 
X"D81", X"D83", X"D86", X"D88", X"D8A", X"D8C", X"D8E", X"D90", 
X"D92", X"D94", X"D97", X"D99", X"D9B", X"D9D", X"D9F", X"DA1", 
X"DA3", X"DA6", X"DA8", X"DAA", X"DAC", X"DAE", X"DB0", X"DB3", 
X"DB5", X"DB7", X"DB9", X"DBB", X"DBD", X"DBF", X"DC1", X"DC4", 
X"DC6", X"DC8", X"DCA", X"DCC", X"DCE", X"DD1", X"DD3", X"DD5", 
X"DD7", X"DD9", X"DDB", X"DDD", X"DE0", X"DE2", X"DE4", X"DE6", 
X"DE8", X"DEA", X"DEC", X"DEE", X"DF1", X"DF3", X"DF5", X"DF7", 
X"DF9", X"DFB", X"DFE", X"E00", X"E02", X"E04", X"E06", X"E08", 
X"E0A", X"E0D", X"E0F", X"E11", X"E13", X"E15", X"E17", X"E19", 
X"E1B", X"E1E", X"E20", X"E22", X"E24", X"E26", X"E28", X"E2B", 
X"E2D", X"E2F", X"E31", X"E33", X"E35", X"E37", X"E3A", X"E3C", 
X"E3E", X"E40", X"E42", X"E44", X"E46", X"E49", X"E4B", X"E4D", 
X"E4F", X"E51", X"E53", X"E55", X"E58", X"E5A", X"E5C", X"E5E", 
X"E60", X"E62", X"E64", X"E67", X"E69", X"E6B", X"E6D", X"E6F", 
X"E71", X"E73", X"E76", X"E78", X"E7A", X"E7C", X"E7E", X"E80", 
X"E82", X"E85", X"E87", X"E89", X"E8B", X"E8D", X"E8F", X"E92", 
X"E94", X"E96", X"E98", X"E9A", X"E9C", X"E9E", X"EA0", X"EA3", 
X"EA5", X"EA7", X"EA9", X"EAB", X"EAD", X"EAF", X"EB2", X"EB4", 
X"EB6", X"EB8", X"EBA", X"EBC", X"EBF", X"EC1", X"EC3", X"EC5", 
X"EC7", X"EC9", X"ECB", X"ECD", X"ED0", X"ED2", X"ED4", X"ED6", 
X"ED8", X"EDA", X"EDC", X"EDF", X"EE1", X"EE3", X"EE5", X"EE7", 
X"EE9", X"EEC", X"EEE", X"EF0", X"EF2", X"EF4", X"EF6", X"EF8", 
X"EFB", X"EFD", X"EFF", X"F01", X"F03", X"F05", X"F07", X"F0A", 
X"F0C", X"F0E", X"F10", X"F12", X"F14", X"F16", X"F19", X"F1B", 
X"F1D", X"F1F", X"F21", X"F23", X"F25", X"F28", X"F2A", X"F2C", 
X"F2E", X"F30", X"F32", X"F34", X"E8B", X"E8D", X"E8F", X"E91", 
X"E93", X"E95", X"E97", X"E9A", X"E9C", X"E9E", X"EA0", X"EA2", 
X"EA4", X"EA7", X"EA9", X"EAB", X"EAD", X"EAF", X"EB1", X"EB3", 
X"EB6", X"EB8", X"EBA", X"EBC", X"EBE", X"EC0", X"EC2", X"EC4", 
X"EC7", X"EC9", X"ECB", X"ECD", X"ECF", X"ED1", X"ED4", X"ED6", 
X"ED8", X"EDA", X"EDC", X"EDE", X"EE0", X"EE3", X"EE5", X"EE7", 
X"EE9", X"EEB", X"EED", X"EEF", X"EF1", X"EF4", X"EF6", X"EF8", 
X"EFA", X"EFC", X"EFE", X"F01", X"F03", X"F05", X"F07", X"F09", 
X"F0B", X"F0D", X"F10", X"F12", X"F14", X"F16", X"F18", X"F1A", 
X"F1C", X"F1F", X"F21", X"F23", X"F25", X"F27", X"F29", X"F2B", 
X"F2E", X"F30", X"F32", X"F34", X"F36", X"F38", X"F3A", X"F3D", 
X"F3F", X"F41", X"F43", X"F45", X"F47", X"F49", X"F4C", X"F4E", 
X"F50", X"F52", X"F54", X"F56", X"F58", X"F5B", X"F5D", X"F5F", 
X"F61", X"F63", X"F65", X"F68", X"F6A", X"F6C", X"F6E", X"F70", 
X"F72", X"F74", X"F76", X"F79", X"F7B", X"F7D", X"F7F", X"F81", 
X"F83", X"F85", X"F88", X"F8A", X"F8C", X"F8E", X"F90", X"F92", 
X"F95", X"F97", X"F99", X"F9B", X"F9D", X"F9F", X"FA1", X"FA3", 
X"FA6", X"FA8", X"FAA", X"FAC", X"FAE", X"FB0", X"FB2", X"FB5", 
X"FB7", X"FB9", X"FBB", X"FBD", X"FBF", X"FC2", X"FC4", X"FC6", 
X"FC8", X"FCA", X"FCC", X"FCE", X"FD0", X"FD3", X"FD5", X"FD7", 
X"FD9", X"FDB", X"FDD", X"FE0", X"FE2", X"FE4", X"FE6", X"FE8", 
X"FEA", X"FEC", X"FEF", X"FF1", X"FF3", X"FF5", X"FF7", X"FF9", 
X"FFB", X"FFD", X"000", X"002", X"004", X"006", X"008", X"00A", 
X"00D", X"00F", X"011", X"013", X"015", X"017", X"019", X"01C", 
X"01E", X"020", X"022", X"024", X"026", X"028", X"02A", X"02D", 
X"02F", X"031", X"033", X"035", X"037", X"03A", X"03C", X"03E", 
X"040", X"042", X"044", X"046", X"049", X"04B", X"04D", X"04F", 
X"051", X"053", X"055", X"057", X"05A", X"05C", X"05E", X"060", 
X"062", X"064", X"067", X"069", X"06B", X"06D", X"06F", X"071", 
X"073", X"076", X"078", X"07A", X"07C", X"07E", X"080", X"082", 
X"085", X"087", X"089", X"08B", X"08D", X"08F", X"091", X"094", 
X"096", X"098", X"09A", X"09C", X"09E", X"0A0", X"0A3", X"0A5", 
X"0A7", X"0A9", X"0AB", X"0AD", X"0AF", X"0B2", X"0B4", X"0B6", 
X"0B8", X"0BA", X"0BC", X"0BE", X"0C1", X"0C3", X"0C5", X"0C7", 
X"0C9", X"0CB", X"0CE", X"0D0", X"0D2", X"0D4", X"0D6", X"0D8", 
X"0DA", X"0DC", X"0DF", X"0E1", X"0E3", X"0E5", X"0E7", X"0E9", 
X"0EB", X"0EE", X"0F0", X"0F2", X"0F4", X"0F6", X"0F8", X"0FB", 
X"0FD", X"0FF", X"101", X"103", X"105", X"107", X"109", X"10C", 
X"10E", X"110", X"112", X"114", X"116", X"118", X"11B", X"11D", 
X"11F", X"121", X"123", X"125", X"128", X"12A", X"12C", X"12E", 
X"130", X"132", X"134", X"137", X"139", X"13B", X"13D", X"13F", 
X"141", X"143", X"146", X"148", X"14A", X"14C", X"14E", X"150", 
X"152", X"155", X"157", X"159", X"15B", X"15D", X"15F", X"161", 
X"164", X"166", X"168", X"16A", X"16C", X"16E", X"170", X"173", 
X"175", X"177", X"179", X"167", X"169", X"16B", X"16D", X"16F", 
X"171", X"173", X"176", X"178", X"17A", X"17C", X"17E", X"180", 
X"183", X"185", X"187", X"189", X"18B", X"18D", X"18F", X"192", 
X"194", X"196", X"198", X"19A", X"19C", X"19E", X"1A0", X"1A3", 
X"1A5", X"1A7", X"1A9", X"1AB", X"1AD", X"1B0", X"1B2", X"1B4", 
X"1B6", X"1B8", X"1BA", X"1BC", X"1BF", X"1C1", X"1C3", X"1C5", 
X"1C7", X"1C9", X"1CB", X"1CD", X"1D0", X"1D2", X"1D4", X"1D6", 
X"1D8", X"1DA", X"1DD", X"1DF", X"1E1", X"1E3", X"1E5", X"1E7", 
X"1E9", X"1EC", X"1EE", X"1F0", X"1F2", X"1F4", X"1F6", X"1F8", 
X"1FB", X"1FD", X"1FF", X"201", X"203", X"205", X"207", X"20A", 
X"20C", X"20E", X"210", X"212", X"214", X"217", X"219", X"21B", 
X"21D", X"21F", X"221", X"223", X"225", X"228", X"22A", X"22C", 
X"22E", X"230", X"232", X"234", X"237", X"239", X"23B", X"23D", 
X"23F", X"241", X"244", X"246", X"248", X"24A", X"24C", X"24E", 
X"250", X"253", X"255", X"257", X"259", X"25B", X"25D", X"25F", 
X"261", X"264", X"266", X"268", X"26A", X"26C", X"26E", X"271", 
X"273", X"275", X"277", X"279", X"27B", X"27D", X"280", X"282", 
X"284", X"286", X"288", X"28A", X"28C", X"28E", X"291", X"293", 
X"295", X"297", X"299", X"29B", X"29E", X"2A0", X"2A2", X"2A4", 
X"2A6", X"2A8", X"2AA", X"2AD", X"2AF", X"2B1", X"2B3", X"2B5", 
X"2B7", X"2B9", X"2BC", X"2BE", X"2C0", X"2C2", X"2C4", X"2C6", 
X"2C8", X"2CB", X"2CD", X"2CF", X"2D1", X"2D3", X"2D5", X"2D8", 
X"2DA", X"2DC", X"2DE", X"2E0", X"2E2", X"2E4", X"2E6", X"2E9", 
X"2EB", X"2ED", X"2EF", X"2F1", X"2F3", X"2F5", X"2F8", X"2FA", 
X"2FC", X"2FE", X"300", X"302", X"305", X"307", X"B0A", X"B0C", 
X"B0E", X"B10", X"B12", X"B14", X"B17", X"B19", X"B1B", X"B1D", 
X"B1F", X"B21", X"B23", X"B26", X"B28", X"B2A", X"B2C", X"B2E", 
X"B30", X"B33", X"B35", X"B37", X"B39", X"B3B", X"B3D", X"B3F", 
X"B41", X"B44", X"B46", X"B48", X"B4A", X"B4C", X"B4E", X"B50", 
X"B53", X"B55", X"B57", X"B59", X"B5B", X"B5D", X"B60", X"B62", 
X"B64", X"B66", X"B68", X"B6A", X"B6C", X"B6E", X"B71", X"B73", 
X"B75", X"B77", X"B79", X"B7B", X"B7E", X"B80", X"B82", X"B84", 
X"B86", X"B88", X"B8A", X"B8D", X"B8F", X"B91", X"B93", X"B95", 
X"B97", X"B99", X"B9B", X"B9E", X"BA0", X"BA2", X"BA4", X"BA6", 
X"BA8", X"BAB", X"BAD", X"BAF", X"BB1", X"BB3", X"BB5", X"BB7", 
X"BBA", X"BBC", X"BBE", X"BC0", X"BC2", X"BC4", X"BC6", X"BC8", 
X"BCB", X"BCD", X"BCF", X"BD1", X"BD3", X"BD5", X"BD8", X"BDA", 
X"BDC", X"BDE", X"BE0", X"BE2", X"BE4", X"BE7", X"BE9", X"BEB", 
X"BED", X"BEF", X"BF1", X"BF3", X"BF6", X"BF8", X"BFA", X"BFC", 
X"BFE", X"C00", X"C02", X"C05", X"C07", X"C09", X"C0B", X"C0D", 
X"C0F", X"C11", X"C14", X"C16", X"C18", X"C1A", X"C1C", X"C1E", 
X"C20", X"C23", X"C25", X"C27", X"C29", X"C2B", X"C2D", X"C2F", 
X"C32", X"C34", X"C36", X"C38", X"C3A", X"C3C", X"C3F", X"C41", 
X"C43", X"C45", X"C47", X"C49", X"C4B", X"C4D", X"C50", X"C52", 
X"C54", X"C56", X"C58", X"C5A", X"C5C", X"C5F", X"C61", X"C63", 
X"C65", X"C67", X"C69", X"C6C", X"C6E", X"C70", X"C72", X"C74", 
X"C76", X"C78", X"C7A", X"C7D", X"C7F", X"C81", X"C83", X"C85", 
X"C87", X"C89", X"C8C", X"C8E", X"C90", X"C92", X"C94", X"C96", 
X"C99", X"C9B", X"C9D", X"C9F", X"CA1", X"CA3", X"CA5", X"CA7", 
X"CAA", X"CAC", X"CAE", X"CB0", X"CB2", X"CB4", X"CB6", X"CB9", 
X"CBB", X"CBD", X"CBF", X"CC1", X"CC3", X"CC6", X"CC8", X"CCA", 
X"CCC", X"CCE", X"CD0", X"CD2", X"CD5", X"CD7", X"CD9", X"CDB", 
X"CDD", X"CDF", X"CE1", X"CE4", X"CE6", X"CE8", X"CEA", X"CEC", 
X"CEE", X"CF0", X"CF3", X"CF5", X"CF7", X"CF9", X"CFB", X"CFD", 
X"D00", X"D02", X"D04", X"D06", X"D08", X"D0A", X"D0C", X"D0E", 
X"D11", X"D13", X"D15", X"D17", X"D19", X"D1B", X"D1D", X"D20", 
X"D22", X"D24", X"D26", X"D28", X"D2A", X"D2D", X"D2F", X"D31", 
X"D33", X"D35", X"D37", X"D39", X"D3B", X"D3E", X"D40", X"D42", 
X"D44", X"D46", X"D48", X"D4A", X"D4D", X"D4F", X"D51", X"CA7", 
X"CA9", X"CAB", X"CAE", X"CB0", X"CB2", X"CB4", X"CB6", X"CB8", 
X"CBA", X"CBD", X"CBF", X"CC1", X"CC3", X"CC5", X"CC7", X"CC9", 
X"CCB", X"CCE", X"CD0", X"CD2", X"CD4", X"CD6", X"CD8", X"CDB", 
X"CDD", X"CDF", X"CE1", X"CE3", X"CE5", X"CE7", X"CEA", X"CEC", 
X"CEE", X"CF0", X"CF2", X"CF4", X"CF6", X"CF9", X"CFB", X"CFD", 
X"CFF", X"D01", X"D03", X"D05", X"D08", X"D0A", X"D0C", X"D0E", 
X"D10", X"D12", X"D15", X"D17", X"D19", X"D1B", X"D1D", X"D1F", 
X"D21", X"D23", X"D26", X"D28", X"D2A", X"D2C", X"D2E", X"D30", 
X"D32", X"D35", X"D37", X"D39", X"D3B", X"D3D", X"D3F", X"D42", 
X"D44", X"D46", X"D48", X"D4A", X"D4C", X"D4E", X"D50", X"D53", 
X"D55", X"D57", X"D59", X"D5B", X"D5D", X"D5F", X"D62", X"D64", 
X"D66", X"D68", X"D6A", X"D6C", X"D6F", X"D71", X"D73", X"D75", 
X"D77", X"D79", X"D7B", X"D7D", X"D80", X"D82", X"D84", X"D86", 
X"D88", X"D8A", X"D8C", X"D8F", X"D91", X"D93", X"D95", X"D97", 
X"D99", X"D9C", X"D9E", X"DA0", X"D8D", X"D90", X"D92", X"D94", 
X"D96", X"D98", X"D9A", X"D9D", X"D9F", X"DA1", X"DA3", X"DA5", 
X"DA7", X"DA9", X"DAC", X"DAE", X"DB0", X"DB2", X"DB4", X"DB6", 
X"DB8", X"DBA", X"DBD", X"DBF", X"DC1", X"DC3", X"DC5", X"DC7", 
X"DCA", X"DCC", X"DCE", X"DD0", X"DD2", X"DD4", X"DD6", X"DD9", 
X"DDB", X"DDD", X"DDF", X"DE1", X"DE3", X"DE5", X"DE7", X"DEA", 
X"DEC", X"DEE", X"DF0", X"DF2", X"DF4", X"DF7", X"DF9", X"DFB", 
X"DFD", X"DFF", X"E01", X"E03", X"E06", X"E08", X"E0A", X"E0C", 
X"E0E", X"E10", X"E12", X"E14", X"E17", X"E19", X"E1B", X"E1D", 
X"E1F", X"E21", X"E24", X"E26", X"E28", X"E2A", X"E2C", X"E2E", 
X"E30", X"E33", X"E35", X"E37", X"E39", X"E3B", X"E3D", X"E3F", 
X"E42", X"E44", X"E46", X"E48", X"E4A", X"E4C", X"E4E", X"E51", 
X"E53", X"E55", X"E57", X"E59", X"E5B", X"E5E", X"E60", X"E62", 
X"E64", X"E66", X"E68", X"E6A", X"E6C", X"E6F", X"E71", X"E73", 
X"E75", X"E77", X"E79", X"E7B", X"E7E", X"E80", X"E82", X"E84", 
X"E86", X"E88", X"E8B", X"E8D", X"E8F", X"E91", X"E93", X"E95", 
X"E97", X"E99", X"E9C", X"E9E", X"EA0", X"EA2", X"EA4", X"EA6", 
X"EA8", X"EAB", X"EAD", X"EAF", X"EB1", X"EB3", X"EB5", X"EB8", 
X"EBA", X"EBC", X"EBE", X"EC0", X"EC2", X"EC4", X"EC6", X"EC9", 
X"ECB", X"ECD", X"ECF", X"ED1", X"ED3", X"ED5", X"ED8", X"EDA", 
X"EDC", X"EDE", X"EE0", X"EE2", X"EE5", X"EE7", X"EE9", X"EEB", 
X"EED", X"EEF", X"EF1", X"EF3", X"EF6", X"EF8", X"EFA", X"EFC", 
X"EFE", X"F00", X"F03", X"F05", X"F07", X"F09", X"F0B", X"F0D", 
X"F0F", X"F12", X"F14", X"F16", X"F18", X"F1A", X"F1C", X"F1E", 
X"F20", X"F23", X"F25", X"F27", X"F29", X"F2B", X"F2D", X"F30", 
X"F32", X"F34", X"F36", X"F38", X"F3A", X"F3C", X"F3F", X"F41", 
X"F43", X"F45", X"F47", X"F49", X"F4B", X"F4D", X"F50", X"F52", 
X"F54", X"F56", X"F58", X"F5A", X"F5D", X"F5F", X"F61", X"F63", 
X"F65", X"F67", X"F69", X"F6C", X"F6E", X"F70", X"F72", X"F74", 
X"F76", X"F78", X"F7A", X"F7D", X"F7F", X"F81", X"F83", X"F85", 
X"F87", X"F8A", X"F8C", X"F8E", X"F90", X"F92", X"F94", X"F96", 
X"F99", X"F9B", X"F9D", X"F9F", X"FA1", X"FA3", X"FA5", X"FA8", 
X"FAA", X"FAC", X"FAE", X"FB0", X"FB2", X"FB4", X"FB7", X"FB9", 
X"FBB", X"FBD", X"FBF", X"FC1", X"FC4", X"FC6", X"FC8", X"FCA", 
X"FCC", X"FCE", X"FD0", X"FD2", X"FD5", X"FD7", X"FD9", X"FDB", 
X"FDD", X"FDF", X"FE1", X"FE4", X"FE6", X"FE8", X"FEA", X"FEC", 
X"FEE", X"FF1", X"FF3", X"FF5", X"FF7", X"FF9", X"FFB", X"FFD", 
X"000", X"002", X"004", X"006", X"008", X"00A", X"00C", X"00E", 
X"011", X"013", X"015", X"017", X"019", X"01B", X"01E", X"020", 
X"022", X"024", X"026", X"028", X"02A", X"02D", X"02F", X"031", 
X"033", X"035", X"037", X"039", X"03B", X"03E", X"040", X"042", 
X"044", X"046", X"048", X"04B", X"04D", X"04F", X"051", X"053", 
X"055", X"057", X"05A", X"05C", X"05E", X"060", X"062", X"064", 
X"066", X"069", X"06B", X"06D", X"06F", X"071", X"073", X"075", 
X"078", X"07A", X"07C", X"07E", X"080", X"082", X"085", X"087", 
X"089", X"08B", X"08D", X"08F", X"091", X"093", X"096", X"098", 
X"09A", X"09C", X"09E", X"0A0", X"0A2", X"0A5", X"0A7", X"0A9", 
X"0AB", X"0AD", X"0AF", X"0B2", X"0B4", X"0B6", X"0B8", X"0BA", 
X"0BC", X"0BE", X"0C0", X"0C3", X"0C5", X"0C7", X"0C9", X"0CB", 
X"0CD", X"0CF", X"0D2", X"0D4", X"0D6", X"0D8", X"0DA", X"0DC", 
X"0DF", X"0E1", X"0E3", X"0E5", X"0E7", X"0E9", X"0EB", X"0ED", 
X"0F0", X"0F2", X"0F4", X"0F6", X"0F8", X"0FA", X"0FC", X"0FF", 
X"101", X"103", X"105", X"107", X"109", X"10C", X"10E", X"110", 
X"112", X"114", X"116", X"118", X"11A", X"11D", X"11F", X"121", 
X"123", X"125", X"127", X"12A", X"12C", X"12E", X"130", X"132", 
X"134", X"136", X"139", X"13B", X"13D", X"13F", X"141", X"143", 
X"145", X"147", X"14A", X"14C", X"14E", X"150", X"152", X"154", 
X"157", X"159", X"15B", X"15D", X"15F", X"161", X"163", X"166", 
X"168", X"16A", X"16C", X"16E", X"170", X"172", X"174", X"177", 
X"179", X"17B", X"17D", X"17F", X"181", X"184", X"186", X"188", 
X"18A", X"18C", X"18E", X"190", X"193", X"195", X"197", X"199", 
X"19B", X"19D", X"19F", X"1A1", X"1A4", X"1A6", X"1A8", X"1AA", 
X"1AC", X"1AE", X"1B1", X"1B3", X"1B5", X"1B7", X"1B9", X"1BB", 
X"1BD", X"1C0", X"1C2", X"1C4", X"1C6", X"1C8", X"1CA", X"1CC", 
X"1CF", X"1D1", X"1D3", X"1D5", X"1D7", X"1D9", X"1DB", X"1DE", 
X"1E0", X"1E2", X"1E4", X"1E6", X"1E8", X"1EB", X"1ED", X"1EF", 
X"1F1", X"1F3", X"1F5", X"1F7", X"1F9", X"1FC", X"1FE", X"200", 
X"202", X"204", X"206", X"208", X"20B", X"20D", X"20F", X"211", 
X"213", X"215", X"218", X"21A", X"21C", X"21E", X"220", X"222", 
X"224", X"226", X"229", X"22B", X"22D", X"22F", X"231", X"233", 
X"235", X"238", X"23A", X"23C", X"23E", X"240", X"242", X"245", 
X"247", X"249", X"24B", X"24D", X"24F", X"251", X"253", X"256", 
X"258", X"25A", X"25C", X"25E", X"260", X"262", X"265", X"267", 
X"269", X"26B", X"26D", X"26F", X"272", X"25F", X"261", X"263", 
X"266", X"268", X"26A", X"26C", X"26E", X"270", X"273", X"275", 
X"277", X"279", X"27B", X"27D", X"27F", X"282", X"284", X"286", 
X"288", X"28A", X"28C", X"28E", X"290", X"293", X"295", X"297", 
X"299", X"29B", X"29D", X"2A0", X"2A2", X"2A4", X"2A6", X"2A8", 
X"2AA", X"2AC", X"2AF", X"2B1", X"2B3", X"2B5", X"2B7", X"2B9", 
X"2BB", X"2BD", X"2C0", X"2C2", X"2C4", X"2C6", X"2C8", X"2CA", 
X"2CD", X"2CF", X"2D1", X"2D3", X"2D5", X"2D7", X"2D9", X"2DC", 
X"2DE", X"2E0", X"2E2", X"2E4", X"2E6", X"2E8", X"2EA", X"2ED", 
X"2EF", X"2F1", X"2F3", X"2F5", X"2F7", X"2FA", X"2FC", X"2FE", 
X"300", X"302", X"304", X"306", X"309", X"30B", X"30D", X"30F", 
X"311", X"313", X"315", X"318", X"31A", X"31C", X"31E", X"320", 
X"322", X"324", X"327", X"329", X"32B", X"32D", X"32F", X"331", 
X"334", X"336", X"338", X"33A", X"33C", X"33E", X"340", X"342", 
X"345", X"347", X"349", X"34B", X"34D", X"34F", X"351", X"354", 
X"356", X"358", X"2AE", X"2B0", X"2B2", X"2B5", X"2B7", X"2B9", 
X"2BB", X"2BD", X"2BF", X"2C1", X"2C4", X"2C6", X"2C8", X"2CA", 
X"2CC", X"2CE", X"2D0", X"2D2", X"2D5", X"2D7", X"2D9", X"2DB", 
X"2DD", X"2DF", X"2E2", X"2E4", X"2E6", X"2E8", X"2EA", X"2EC", 
X"2EE", X"2F1", X"2F3", X"2F5", X"2F7", X"2F9", X"2FB", X"2FD", 
X"2FF", X"302", X"304", X"306", X"308", X"30A", X"30C", X"30F", 
X"311", X"313", X"315", X"317", X"319", X"31B", X"31E", X"320", 
X"322", X"324", X"326", X"328", X"32A", X"32D", X"32F", X"331", 
X"333", X"335", X"337", X"339", X"33C", X"33E", X"340", X"342", 
X"344", X"346", X"349", X"34B", X"34D", X"34F", X"351", X"353", 
X"355", X"358", X"35A", X"35C", X"35E", X"360", X"362", X"364", 
X"366", X"369", X"36B", X"36D", X"36F", X"371", X"373", X"376", 
X"378", X"37A", X"37C", X"37E", X"380", X"382", X"385", X"387", 
X"389", X"38B", X"38D", X"38F", X"391", X"393", X"396", X"398", 
X"39A", X"39C", X"39E", X"3A0", X"3A3", X"3A5", X"3A7", X"3A9", 
X"3AB", X"3AD", X"3AF", X"3B2", X"3B4", X"3B6", X"3B8", X"3BA", 
X"3BC", X"3BE", X"3C0", X"3C3", X"3C5", X"3C7", X"3C9", X"3CB", 
X"3CD", X"3D0", X"3D2", X"3D4", X"3D6", X"3D8", X"3DA", X"3DC", 
X"3DF", X"3E1", X"3E3", X"3E5", X"3E7", X"3E9", X"3EB", X"3EE", 
X"3F0", X"3F2", X"3F4", X"3F6", X"3F8", X"3FA", X"3FD", X"3FF", 
X"401", X"403", X"405", X"407", X"409", X"40C", X"40E", X"410", 
X"412", X"414", X"416", X"418", X"41B", X"41D", X"41F", X"421", 
X"423", X"425", X"427", X"42A", X"42C", X"42E", X"430", X"432", 
X"434", X"437", X"439", X"43B", X"43D", X"43F", X"441", X"443", 
X"445", X"448", X"44A", X"44C", X"44E", X"450", X"452", X"454", 
X"457", X"459", X"45B", X"45D", X"45F", X"461", X"464", X"466", 
X"468", X"46A", X"46C", X"46E", X"470", X"472", X"475", X"477", 
X"479", X"47B", X"47D", X"47F", X"481", X"484", X"486", X"488", 
X"48A", X"48C", X"48E", X"491", X"493", X"495", X"497", X"499", 
X"49B", X"49D", X"49F", X"4A2", X"4A4", X"4A6", X"4A8", X"4AA", 
X"4AC", X"4AF", X"4B1", X"4B3", X"4B5", X"4B7", X"4B9", X"4BB", 
X"4BE", X"4C0", X"4C2", X"4C4", X"4C6", X"4C8", X"4CA", X"4CC", 
X"4CF", X"4D1", X"4D3", X"4D5", X"4D7", X"4D9", X"4DC", X"4DE", 
X"4E0", X"4E2", X"4E4", X"4E6", X"4E8", X"4EB", X"4ED", X"4EF", 
X"4F1", X"4F3", X"4F5", X"CF8", X"CFA", X"CFD", X"CFF", X"D01", 
X"D03", X"D05", X"D07", X"D0A", X"D0C", X"D0E", X"D10", X"D12", 
X"D14", X"D16", X"D19", X"D1B", X"D1D", X"D1F", X"D21", X"D23", 
X"D25", X"D27", X"D2A", X"D2C", X"D2E", X"D30", X"D32", X"D34", 
X"D37", X"D39", X"D3B", X"D3D", X"D3F", X"D41", X"D43", X"D46", 
X"D48", X"D4A", X"D4C", X"D4E", X"D50", X"D52", X"D55", X"D57", 
X"D59", X"D5B", X"D5D", X"D5F", X"D61", X"D64", X"D66", X"D68", 
X"D6A", X"D6C", X"D6E", X"D71", X"D73", X"D75", X"D77", X"D79", 
X"D7B", X"D7D", X"D7F", X"D82", X"D84", X"D86", X"D88", X"D8A", 
X"D8C", X"D8E", X"D91", X"D93", X"D95", X"D97", X"D99", X"D9B", 
X"D9E", X"DA0", X"DA2", X"DA4", X"DA6", X"DA8", X"DAA", X"DAC", 
X"DAF", X"DB1", X"DB3", X"DB5", X"DB7", X"DB9", X"DBB", X"DBE", 
X"DC0", X"DC2", X"DC4", X"DC6", X"DC8", X"DCB", X"DCD", X"DCF", 
X"DD1", X"DD3", X"DD5", X"DD7", X"DDA", X"DDC", X"DDE", X"DE0", 
X"DE2", X"DE4", X"DE6", X"DE8", X"DEB", X"DED", X"DEF", X"DF1", 
X"DF3", X"DF5", X"DF8", X"DFA", X"DFC", X"DFE", X"E00", X"E02", 
X"E04", X"E07", X"E09", X"E0B", X"E0D", X"E0F", X"E11", X"E13", 
X"E16", X"E18", X"E1A", X"E1C", X"E1E", X"E20", X"E22", X"E25", 
X"E27", X"E29", X"E2B", X"E2D", X"E2F", X"E32", X"E34", X"E36", 
X"E38", X"E3A", X"E3C", X"E3E", X"E40", X"E43", X"E45", X"E47", 
X"E49", X"E4B", X"E4D", X"E4F", X"E52", X"E54", X"E56", X"E58", 
X"E5A", X"E5C", X"E5F", X"E61", X"E63", X"E65", X"E67", X"E69", 
X"E6B", X"E6D", X"E70", X"E72", X"E74", X"E76", X"E78", X"E7A", 
X"E7C", X"E7F", X"E81", X"E83", X"E85", X"E87", X"E89", X"E8C", 
X"E8E", X"E90", X"E92", X"E94", X"E96", X"E98", X"E86", X"E88", 
X"E8A", X"E8C", X"E8F", X"E91", X"E93", X"E95", X"E97", X"E99", 
X"E9B", X"E9E", X"EA0", X"EA2", X"EA4", X"EA6", X"EA8", X"EAA", 
X"EAD", X"EAF", X"EB1", X"EB3", X"EB5", X"EB7", X"EB9", X"EBC", 
X"EBE", X"EC0", X"EC2", X"EC4", X"EC6", X"EC8", X"ECB", X"ECD", 
X"ECF", X"ED1", X"ED3", X"ED5", X"ED7", X"EDA", X"EDC", X"EDE", 
X"EE0", X"EE2", X"EE4", X"EE7", X"EE9", X"EEB", X"EED", X"EEF", 
X"EF1", X"EF3", X"EF6", X"EF8", X"EFA", X"EFC", X"EFE", X"F00", 
X"F02", X"F04", X"F07", X"F09", X"F0B", X"F0D", X"F0F", X"F11", 
X"F14", X"F16", X"F18", X"F1A", X"F1C", X"F1E", X"F20", X"F23", 
X"F25", X"F27", X"F29", X"F2B", X"F2D", X"F2F", X"F31", X"F34", 
X"F36", X"F38", X"F3A", X"F3C", X"F3E", X"F41", X"F43", X"F45", 
X"F47", X"F49", X"F4B", X"F4D", X"F50", X"F52", X"F54", X"F56", 
X"F58", X"F5A", X"F5C", X"F5F", X"F61", X"F63", X"F65", X"F67", 
X"F69", X"F6B", X"F6E", X"F70", X"F72", X"F74", X"F76", X"F78", 
X"F7A", X"F7D", X"F7F", X"F81", X"F83", X"F85", X"F87", X"F89", 
X"F8C", X"F8E", X"F90", X"F92", X"F94", X"F96", X"F98", X"F9B", 
X"F9D", X"F9F", X"FA1", X"FA3", X"FA5", X"FA8", X"FAA", X"FAC", 
X"FAE", X"FB0", X"FB2", X"FB4", X"FB6", X"FB9", X"FBB", X"FBD", 
X"FBF", X"FC1", X"FC3", X"FC5", X"FC8", X"FCA", X"FCC", X"FCE", 
X"FD0", X"FD2", X"FD5", X"FD7", X"FD9", X"FDB", X"FDD", X"FDF", 
X"FE1", X"FE3", X"FE6", X"FE8", X"FEA", X"FEC", X"FEE", X"FF0", 
X"FF2", X"FF5", X"FF7", X"FF9", X"FFB", X"FFD", X"FFF", X"002", 
X"004", X"006", X"008", X"00A", X"00C", X"00E", X"010", X"013", 
X"015", X"017", X"019", X"01B", X"01D", X"01F", X"022", X"024", 
X"026", X"028", X"02A", X"02C", X"02F", X"031", X"033", X"035", 
X"037", X"039", X"03B", X"03D", X"040", X"042", X"044", X"046", 
X"048", X"04A", X"04D", X"04F", X"051", X"053", X"055", X"057", 
X"059", X"05C", X"05E", X"060", X"062", X"064", X"066", X"068", 
X"06A", X"06D", X"06F", X"071", X"073", X"075", X"077", X"07A", 
X"07C", X"07E", X"080", X"082", X"084", X"086", X"089", X"08B", 
X"08D", X"08F", X"091", X"093", X"095", X"097", X"09A", X"09C", 
X"09E", X"0A0", X"0A2", X"0A4", X"0A7", X"0A9", X"0AB", X"0AD", 
X"0AF", X"0B1", X"0B3", X"0B6", X"0B8", X"0BA", X"0BC", X"0BE", 
X"0C0", X"0C2", X"0C5", X"0C7", X"0C9", X"0CB", X"0CD", X"0CF", 
X"0D1", X"0D4", X"0D6", X"0D8", X"0DA", X"0DC", X"0DE", X"0E0", 
X"0E3", X"0E5", X"0E7", X"0E9", X"0EB", X"0ED", X"0EF", X"0F2", 
X"0F4", X"0F6", X"0F8", X"0FA", X"0FC", X"0FE", X"101", X"103", 
X"105", X"107", X"109", X"10B", X"10E", X"110", X"112", X"114", 
X"116", X"118", X"11A", X"11C", X"11F", X"121", X"123", X"125", 
X"127", X"129", X"12B", X"12E", X"130", X"132", X"134", X"136", 
X"138", X"13B", X"13D", X"13F", X"141", X"143", X"145", X"147", 
X"149", X"14C", X"14E", X"150", X"152", X"154", X"156", X"158", 
X"15B", X"15D", X"15F", X"161", X"163", X"165", X"168", X"16A", 
X"16C", X"16E", X"170", X"172", X"174", X"0CB", X"0CD", X"0CF", 
X"0D1", X"0D3", X"0D5", X"0D7", X"0DA", X"0DC", X"0DE", X"0E0", 
X"0E2", X"0E4", X"0E6", X"0E9", X"0EB", X"0ED", X"0EF", X"0F1", 
X"0F3", X"0F5", X"0F8", X"0FA", X"0FC", X"0FE", X"100", X"102", 
X"104", X"107", X"109", X"10B", X"10D", X"10F", X"111", X"113", 
X"116", X"118", X"11A", X"11C", X"11E", X"120", X"123", X"125", 
X"127", X"129", X"12B", X"12D", X"12F", X"132", X"134", X"136", 
X"138", X"13A", X"13C", X"13E", X"140", X"143", X"145", X"147", 
X"149", X"14B", X"14D", X"150", X"152", X"154", X"156", X"158", 
X"15A", X"15C", X"15F", X"161", X"163", X"165", X"167", X"169", 
X"16B", X"16D", X"170", X"172", X"174", X"176", X"178", X"17A", 
X"17D", X"17F", X"181", X"183", X"185", X"187", X"189", X"18C", 
X"18E", X"190", X"192", X"194", X"196", X"198", X"19B", X"19D", 
X"19F", X"1A1", X"1A3", X"1A5", X"1A7", X"1AA", X"1AC", X"1AE", 
X"1B0", X"1B2", X"1B4", X"1B6", X"1B9", X"1BB", X"1BD", X"1BF", 
X"1C1", X"1C3", X"1C5", X"1C8", X"1CA", X"1CC", X"1CE", X"1D0", 
X"1D2", X"1D4", X"1D7", X"1D9", X"1DB", X"1DD", X"1DF", X"1E1", 
X"1E4", X"1E6", X"1E8", X"1EA", X"1EC", X"1EE", X"1F0", X"1F2", 
X"1F5", X"1F7", X"1F9", X"1FB", X"1FD", X"1FF", X"201", X"204", 
X"206", X"208", X"20A", X"20C", X"20E", X"211", X"213", X"215", 
X"217", X"219", X"21B", X"21D", X"21F", X"222", X"224", X"226", 
X"228", X"22A", X"22C", X"22E", X"231", X"233", X"235", X"237", 
X"239", X"23B", X"23E", X"240", X"242", X"244", X"246", X"248", 
X"24A", X"24C", X"24F", X"251", X"253", X"255", X"257", X"259", 
X"25C", X"25E", X"260", X"262", X"264", X"266", X"268", X"26B", 
X"26D", X"26F", X"271", X"273", X"275", X"277", X"279", X"27C", 
X"27E", X"280", X"282", X"284", X"286", X"289", X"28B", X"28D", 
X"28F", X"291", X"293", X"295", X"298", X"29A", X"29C", X"29E", 
X"2A0", X"2A2", X"2A4", X"2A6", X"2A9", X"2AB", X"2AD", X"2AF", 
X"2B1", X"2B3", X"2B6", X"2B8", X"2BA", X"2BC", X"2BE", X"2AC", 
X"2AE", X"2B0", X"2B2", X"2B4", X"2B6", X"2B9", X"2BB", X"2BD", 
X"2BF", X"2C1", X"2C3", X"2C6", X"2C8", X"2CA", X"2CC", X"2CE", 
X"2D0", X"2D2", X"2D5", X"2D7", X"2D9", X"2DB", X"2DD", X"2DF", 
X"2E1", X"2E3", X"2E6", X"2E8", X"2EA", X"2EC", X"2EE", X"2F0", 
X"2F3", X"2F5", X"2F7", X"2F9", X"2FB", X"2FD", X"2FF", X"302", 
X"304", X"306", X"308", X"30A", X"30C", X"30E", X"311", X"313", 
X"315", X"317", X"319", X"31B", X"31D", X"320", X"322", X"324", 
X"326", X"328", X"32A", X"32D", X"32F", X"331", X"333", X"335", 
X"337", X"339", X"33B", X"33E", X"340", X"342", X"344", X"346", 
X"348", X"34A", X"34D", X"34F", X"351", X"353", X"355", X"357", 
X"35A", X"35C", X"35E", X"360", X"362", X"364", X"366", X"368", 
X"36B", X"36D", X"36F", X"371", X"373", X"375", X"377", X"37A", 
X"37C", X"37E", X"380", X"382", X"384", X"387", X"389", X"38B", 
X"38D", X"38F", X"391", X"393", X"395", X"398", X"39A", X"39C", 
X"39E", X"3A0", X"3A2", X"3A4", X"3A7", X"3A9", X"3AB", X"3AD", 
X"3AF", X"3B1", X"3B4", X"3B6", X"3B8", X"3BA", X"3BC", X"3BE", 
X"3C0", X"3C2", X"3C5", X"3C7", X"3C9", X"3CB", X"3CD", X"3CF", 
X"3D2", X"3D4", X"3D6", X"3D8", X"3DA", X"3DC", X"3DE", X"3E1", 
X"3E3", X"3E5", X"3E7", X"3E9", X"3EB", X"3ED", X"3EF", X"3F2", 
X"3F4", X"3F6", X"3F8", X"3FA", X"3FC", X"3FF", X"401", X"403", 
X"405", X"407", X"409", X"40B", X"40E", X"410", X"412", X"414", 
X"416", X"418", X"41A", X"41C", X"41F", X"421", X"423", X"425", 
X"427", X"429", X"42C", X"42E", X"430", X"432", X"434", X"436", 
X"438", X"43B", X"43D", X"43F", X"441", X"443", X"445", X"447", 
X"449", X"44C", X"44E", X"450", X"452", X"454", X"456", X"459", 
X"45B", X"45D", X"45F", X"461", X"463", X"465", X"468", X"46A", 
X"46C", X"46E", X"470", X"472", X"474", X"477", X"479", X"47B", 
X"47D", X"47F", X"481", X"483", X"486", X"488", X"48A", X"48C", 
X"48E", X"490", X"493", X"495", X"497", X"499", X"49B", X"49D", 
X"49F", X"4A1", X"4A4", X"4A6", X"4A8", X"4AA", X"4AC", X"4AE", 
X"4B0", X"4B3", X"4B5", X"4B7", X"4B9", X"4BB", X"4BD", X"4C0", 
X"4C2", X"4C4", X"4C6", X"4C8", X"4CA", X"4CC", X"4CF", X"4D1", 
X"4D3", X"4D5", X"4D7", X"4D9", X"4DB", X"4DD", X"4E0", X"4E2", 
X"4E4", X"4E6", X"4E8", X"4EA", X"4ED", X"4EF", X"4F1", X"4F3", 
X"4F5", X"4F7", X"4F9", X"4FC", X"4FE", X"500", X"502", X"504", 
X"506", X"508", X"50A", X"50D", X"50F", X"511", X"513", X"515", 
X"517", X"51A", X"51C", X"51E", X"520", X"522", X"524", X"526", 
X"529", X"52B", X"52D", X"52F", X"531", X"533", X"535", X"538", 
X"53A", X"53C", X"53E", X"540", X"542", X"544", X"547", X"549", 
X"54B", X"54D", X"54F", X"551", X"554", X"556", X"558", X"55A", 
X"55C", X"55E", X"560", X"562", X"565", X"567", X"569", X"56B", 
X"56D", X"56F", X"571", X"574", X"576", X"578", X"57A", X"57C", 
X"57E", X"581", X"583", X"585", X"587", X"589", X"58B", X"58D", 
X"58F", X"592", X"594", X"596", X"598", X"59A", X"59C", X"59E", 
X"5A1", X"5A3", X"5A5", X"5A7", X"5A9", X"5AB", X"5AE", X"5B0", 
X"5B2", X"5B4", X"5B6", X"5B8", X"5BA", X"5BC", X"5BF", X"5C1", 
X"5C3", X"5C5", X"5C7", X"5C9", X"5CB", X"5CE", X"5D0", X"5D2", 
X"5D4", X"5D6", X"5D8", X"5DB", X"5DD", X"5DF", X"5E1", X"5E3", 
X"5E5", X"5E7", X"5E9", X"5EC", X"5EE", X"5F0", X"5F2", X"5F4", 
X"5F6", X"5F9", X"5FB", X"5FD", X"5FF", X"601", X"603", X"605", 
X"608", X"60A", X"60C", X"60E", X"610", X"612", X"614", X"616", 
X"619", X"61B", X"61D", X"61F", X"621", X"623", X"626", X"628", 
X"62A", X"62C", X"62E", X"630", X"632", X"635", X"637", X"639", 
X"63B", X"63D", X"63F", X"641", X"643", X"646", X"648", X"64A", 
X"64C", X"64E", X"650", X"653", X"655", X"657", X"659", X"65B", 
X"65D", X"65F", X"662", X"664", X"666", X"668", X"66A", X"66C", 
X"66E", X"671", X"673", X"675", X"677", X"679", X"67B", X"67D", 
X"680", X"682", X"684", X"686", X"688", X"68A", X"68C", X"68F", 
X"691", X"693", X"695", X"697", X"699", X"69B", X"69E", X"6A0", 
X"6A2", X"6A4", X"6A6", X"6A8", X"6AA", X"6AD", X"6AF", X"6B1", 
X"6B3", X"6B5", X"6B7", X"6BA", X"6BC", X"6BE", X"6C0", X"6C2", 
X"6C4", X"6C6", X"6C8", X"6CB", X"6CD", X"6CF", X"6D1", X"6D3", 
X"6D5", X"6D7", X"6DA", X"6DC", X"6DE", X"6E0", X"6E2", X"6E4", 
X"6E7", X"6E9", X"6EB", X"6ED", X"6EF", X"6F1", X"6F3", X"6F5", 
X"6F8", X"6FA", X"6FC", X"6FE", X"700", X"702", X"704", X"707", 
X"709", X"70B", X"70D", X"70F", X"711", X"714", X"716", X"718", 
X"71A", X"71C", X"71E", X"720", X"722", X"725", X"727", X"729", 
X"72B", X"72D", X"72F", X"732", X"734", X"736", X"738", X"73A", 
X"73C", X"73E", X"741", X"743", X"745", X"747", X"749", X"74B", 
X"74D", X"74F", X"752", X"754", X"756", X"758", X"75A", X"75C", 
X"75F", X"761", X"763", X"765", X"767", X"769", X"76B", X"76E", 
X"770", X"772", X"774", X"776", X"778", X"77B", X"77D", X"77F", 
X"781", X"783", X"785", X"787", X"789", X"78C", X"78E", X"790"
);

signal data : std_logic_vector(31 downto 0);
signal unsignedIndex : unsigned(11 downto 0) := X"000";

begin

rom_select: process (clk, en)
begin
	if (rising_edge(clk)) then
    if (en = '1') then
		unsignedIndex <= unsigned(address_reg);
		data <= (SIN_ROM(to_integer(unsignedIndex)) & x"00000");
		sin_out <= std_logic_vector(shift_right(signed(data), 20));
    end if;
  end if;
end process rom_select;

end rtl;
