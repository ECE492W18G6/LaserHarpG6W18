  --------------------------------------------------------------------------------------------------------------------------
-- Original Authors : Simon Doherty, Eric Lunty, Kyle Brooks, Peter Roland						--
-- Date created: N/A 													--
--															--
-- Additional Authors : Randi Derbyshire, Adam Narten, Oliver Rarog, Celeste Chiasson					--
-- Date edited: March 26, 2018											--
--															--
-- This program takes a value from the synthesizer.vhd file and runs it through the 12-bit ROM to find the 	 	--
-- respective sine wave value. 												--
--------------------------------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use IEEE.STD_LOGIC_SIGNED.all;
use ieee.numeric_std.all;               -- Needed for shifts

entity ClarinetSin_lut is

port (
	clk      : in  std_logic;
	en       : in  std_logic;
	
	--Address input
	address_reg : in std_logic_vector(11 downto 0); 
	
	--Sine value output
	sin_out  : out std_logic_vector(31 downto 0)
	);
end entity;


architecture rtl of ClarinetSin_lut is


type rom_type is array (0 to 4095) of std_logic_vector (11 downto 0);

constant SIN_ROM : rom_type :=

(
X"000", X"00D", X"01A", X"026", X"033", X"040", X"04D", X"059", 
X"066", X"073", X"080", X"08C", X"099", X"0A6", X"0B3", X"0BF", 
X"0CC", X"0D8", X"0E5", X"0F2", X"0FE", X"10B", X"118", X"124", 
X"130", X"13D", X"149", X"156", X"162", X"16E", X"17B", X"187", 
X"194", X"19F", X"1AC", X"1B8", X"1C4", X"1D0", X"1DC", X"1E8", 
X"1F4", X"1FF", X"20B", X"218", X"224", X"22E", X"23A", X"246", 
X"252", X"25E", X"268", X"274", X"27F", X"28B", X"295", X"2A1", 
X"2AC", X"2B7", X"2C2", X"2CD", X"2D8", X"2E3", X"2EE", X"2F8", 
X"303", X"30D", X"318", X"322", X"32C", X"337", X"341", X"34B", 
X"355", X"35F", X"369", X"372", X"37C", X"386", X"390", X"39A", 
X"3A3", X"3AC", X"3B6", X"3BF", X"3C8", X"3D1", X"3DA", X"3E3", 
X"3EC", X"3F5", X"3FE", X"406", X"40F", X"417", X"420", X"428", 
X"430", X"438", X"440", X"448", X"450", X"458", X"460", X"467", 
X"46F", X"476", X"47E", X"485", X"48C", X"494", X"49A", X"4A1", 
X"4A8", X"4AF", X"4B6", X"4BC", X"4C3", X"4CA", X"4D0", X"4D6", 
X"4DC", X"4E3", X"4E9", X"4EE", X"4F4", X"4FA", X"500", X"505", 
X"50B", X"511", X"516", X"51B", X"520", X"525", X"52B", X"52F", 
X"534", X"539", X"53E", X"543", X"547", X"54B", X"550", X"554", 
X"558", X"55C", X"561", X"565", X"568", X"56C", X"570", X"574", 
X"577", X"57B", X"57E", X"582", X"585", X"588", X"58B", X"58E", 
X"591", X"594", X"597", X"59A", X"59D", X"59F", X"5A2", X"5A4", 
X"5A7", X"5A9", X"5AB", X"5AE", X"5B0", X"5B2", X"5B4", X"5B6", 
X"5B8", X"5BA", X"5BB", X"5BD", X"5BF", X"5C0", X"5C2", X"5C3", 
X"5C5", X"5C6", X"5C7", X"5C9", X"5CA", X"5CB", X"5CC", X"5CD", 
X"5CE", X"5CF", X"5D0", X"5D0", X"5D1", X"5D2", X"5D2", X"5D3", 
X"5D4", X"5D4", X"5D4", X"5D5", X"5D5", X"5D5", X"5D6", X"5D6", 
X"5D6", X"5D6", X"5D6", X"5D6", X"5D6", X"5D6", X"5D6", X"5D6", 
X"5D6", X"5D6", X"5D6", X"5D5", X"5D5", X"5D5", X"5D4", X"5D4", 
X"5D3", X"5D3", X"5D2", X"5D2", X"5D1", X"5D1", X"5D0", X"5CF", 
X"5CF", X"5CE", X"5CD", X"5CC", X"5CC", X"5CB", X"5CA", X"5C9", 
X"5C8", X"5C7", X"5C6", X"5C5", X"5C4", X"5C3", X"5C2", X"5C1", 
X"5C0", X"5BF", X"5BE", X"5BD", X"5BC", X"5BB", X"5BA", X"5B8", 
X"5B7", X"5B6", X"5B5", X"5B3", X"5B2", X"5B1", X"5B0", X"5AE", 
X"5AD", X"5AC", X"5AB", X"5A9", X"5A8", X"5A7", X"5A5", X"5A4", 
X"5A2", X"5A1", X"5A0", X"59E", X"59D", X"59C", X"59A", X"599", 
X"597", X"596", X"595", X"593", X"592", X"590", X"58F", X"58D", 
X"58C", X"58A", X"589", X"588", X"586", X"585", X"583", X"582", 
X"580", X"57F", X"57E", X"57C", X"57B", X"579", X"578", X"576", 
X"575", X"573", X"572", X"571", X"56F", X"56E", X"56C", X"56B", 
X"569", X"568", X"567", X"565", X"564", X"562", X"561", X"55F", 
X"55E", X"55D", X"55B", X"55A", X"559", X"557", X"556", X"554", 
X"553", X"552", X"550", X"54F", X"54E", X"54C", X"54B", X"54A", 
X"548", X"547", X"546", X"544", X"543", X"542", X"541", X"53F", 
X"53E", X"53D", X"53B", X"53A", X"539", X"538", X"536", X"535", 
X"534", X"533", X"531", X"530", X"52F", X"52E", X"52C", X"52B", 
X"52A", X"529", X"528", X"526", X"525", X"524", X"523", X"522", 
X"520", X"51F", X"51E", X"51D", X"51C", X"51B", X"519", X"518", 
X"517", X"516", X"515", X"514", X"513", X"512", X"510", X"50F", 
X"50E", X"50D", X"50C", X"50B", X"50A", X"509", X"507", X"506", 
X"505", X"504", X"503", X"502", X"501", X"500", X"4FF", X"4FE", 
X"4FD", X"4FC", X"4FA", X"4F9", X"4F8", X"4F7", X"4F6", X"4F5", 
X"4F4", X"4F3", X"4F2", X"4F1", X"4F0", X"4EF", X"4EE", X"4ED", 
X"4EC", X"4EB", X"4EA", X"4E9", X"4E7", X"4E6", X"4E5", X"4E4", 
X"4E3", X"4E2", X"4E1", X"4E0", X"4DF", X"4DE", X"4DD", X"4DC", 
X"4DB", X"4DA", X"4D9", X"4D8", X"4D7", X"4D6", X"4D5", X"4D4", 
X"4D3", X"4D2", X"4D1", X"4D0", X"4CF", X"4CE", X"4CD", X"4CC", 
X"4CB", X"4CA", X"4C9", X"4C8", X"4C7", X"4C6", X"4C5", X"4C4", 
X"4C3", X"4C2", X"4C1", X"4C0", X"4BF", X"4BE", X"4BD", X"4BC", 
X"4BB", X"4BA", X"4B9", X"4B8", X"4B7", X"4B6", X"4B5", X"4B4", 
X"4B3", X"4B2", X"4B1", X"4B0", X"4AF", X"4AE", X"4AD", X"4AC", 
X"4AB", X"4AA", X"4A9", X"4A8", X"4A7", X"4A6", X"4A5", X"4A4", 
X"4A3", X"4A2", X"4A2", X"4A1", X"4A0", X"49F", X"49E", X"49D", 
X"49C", X"49B", X"49A", X"499", X"498", X"497", X"496", X"495", 
X"494", X"493", X"492", X"491", X"490", X"490", X"48F", X"48E", 
X"48D", X"48C", X"48B", X"48A", X"489", X"488", X"487", X"486", 
X"485", X"484", X"483", X"482", X"481", X"481", X"480", X"47F", 
X"47E", X"47D", X"47C", X"47B", X"47A", X"479", X"478", X"477", 
X"476", X"475", X"474", X"473", X"472", X"471", X"470", X"46F", 
X"46E", X"46D", X"46C", X"46C", X"46B", X"46A", X"469", X"468", 
X"467", X"466", X"465", X"464", X"463", X"462", X"461", X"460", 
X"45F", X"45D", X"45C", X"45B", X"45A", X"459", X"458", X"457", 
X"456", X"455", X"454", X"453", X"452", X"451", X"44F", X"44E", 
X"44D", X"44C", X"44B", X"44A", X"448", X"447", X"446", X"445", 
X"444", X"443", X"441", X"440", X"43F", X"43D", X"43C", X"43B", 
X"43A", X"438", X"437", X"436", X"434", X"433", X"431", X"430", 
X"42F", X"42D", X"42C", X"42A", X"429", X"427", X"426", X"424", 
X"423", X"421", X"41F", X"41E", X"41C", X"41B", X"419", X"417", 
X"416", X"414", X"412", X"410", X"40F", X"40D", X"40B", X"409", 
X"407", X"405", X"403", X"401", X"400", X"3FE", X"3FC", X"3FA", 
X"3F8", X"3F6", X"3F3", X"3F1", X"3EF", X"3ED", X"3EB", X"3E9", 
X"3E6", X"3E4", X"3E2", X"3DF", X"3DD", X"3DB", X"3D8", X"3D6", 
X"3D3", X"3D1", X"3CF", X"3CC", X"3C9", X"3C7", X"3C4", X"3C2", 
X"3BF", X"3BC", X"3BA", X"3B7", X"3B4", X"3B1", X"3AF", X"3AC", 
X"3A9", X"3A6", X"3A3", X"3A0", X"39D", X"39A", X"397", X"394", 
X"390", X"38D", X"38A", X"387", X"384", X"380", X"37D", X"379", 
X"376", X"373", X"36F", X"36C", X"368", X"365", X"361", X"35E", 
X"35A", X"356", X"353", X"34F", X"34B", X"347", X"344", X"340", 
X"33C", X"338", X"334", X"330", X"32C", X"328", X"324", X"320", 
X"31C", X"318", X"313", X"30F", X"30B", X"306", X"302", X"2FE", 
X"2FA", X"2F5", X"2F1", X"2EC", X"2E8", X"2E3", X"2DF", X"2DA", 
X"2D6", X"2D1", X"2CD", X"2C8", X"2C3", X"2BE", X"2BA", X"2B5", 
X"2B0", X"2AB", X"2A6", X"2A2", X"29D", X"298", X"293", X"28E", 
X"289", X"284", X"27F", X"27A", X"275", X"270", X"26A", X"265", 
X"260", X"25B", X"256", X"250", X"24B", X"246", X"241", X"23B", 
X"236", X"231", X"22B", X"226", X"220", X"21B", X"216", X"210", 
X"20B", X"206", X"200", X"1FA", X"1F5", X"1F0", X"1EA", X"1E4", 
X"1DF", X"1D9", X"1D4", X"1CE", X"1C8", X"1C3", X"1BE", X"1B8", 
X"1B2", X"1AC", X"1A7", X"1A1", X"19C", X"196", X"190", X"18B", 
X"185", X"17F", X"179", X"174", X"16E", X"168", X"163", X"15D", 
X"158", X"152", X"14C", X"147", X"141", X"13B", X"135", X"12F", 
X"12A", X"124", X"11F", X"119", X"114", X"10E", X"108", X"102", 
X"0FD", X"0F7", X"0F2", X"0EC", X"0E7", X"0E1", X"0DB", X"0D6", 
X"0D0", X"0CB", X"0C5", X"0C0", X"0BA", X"0B5", X"0AF", X"0AA", 
X"0A4", X"09F", X"099", X"094", X"08E", X"089", X"084", X"07F", 
X"079", X"074", X"06F", X"069", X"064", X"05F", X"05A", X"055", 
X"04F", X"04A", X"045", X"040", X"03B", X"036", X"031", X"02C", 
X"027", X"022", X"01D", X"018", X"013", X"00E", X"009", X"005", 
X"000", X"FFB", X"FF6", X"FF1", X"FED", X"FE8", X"FE4", X"FDF", 
X"FDB", X"FD6", X"FD1", X"FCD", X"FC9", X"FC4", X"FC0", X"FBB", 
X"FB7", X"FB3", X"FAE", X"FAA", X"FA6", X"FA2", X"F9E", X"F99", 
X"F95", X"F91", X"F8D", X"F89", X"F85", X"F82", X"F7E", X"F7A", 
X"F76", X"F72", X"F6E", X"F6A", X"F67", X"F63", X"F5F", X"F5C", 
X"F58", X"F54", X"F51", X"F4E", X"F4A", X"F47", X"F43", X"F40", 
X"F3D", X"F39", X"F36", X"F33", X"F30", X"F2C", X"F29", X"F26", 
X"F23", X"F20", X"F1D", X"F1A", X"F17", X"F14", X"F11", X"F0F", 
X"F0C", X"F09", X"F06", X"F03", X"F01", X"EFE", X"EFC", X"EF9", 
X"EF7", X"EF4", X"EF2", X"EEF", X"EED", X"EEA", X"EE8", X"EE6", 
X"EE3", X"EE1", X"EDF", X"EDD", X"EDA", X"ED8", X"ED6", X"ED4", 
X"ED2", X"ED0", X"ECE", X"ECC", X"ECA", X"EC8", X"EC6", X"EC4", 
X"EC3", X"EC1", X"EBF", X"EBD", X"EBC", X"EBA", X"EB8", X"EB7", 
X"EB5", X"EB4", X"EB2", X"EB1", X"EAF", X"EAE", X"EAC", X"EAB", 
X"EA9", X"EA8", X"EA7", X"EA6", X"EA4", X"EA3", X"EA2", X"EA1", 
X"EA0", X"E9E", X"E9D", X"E9C", X"E9B", X"E9A", X"E99", X"E98", 
X"E97", X"E96", X"E95", X"E94", X"E94", X"E93", X"E92", X"E91", 
X"E91", X"E90", X"E8F", X"E8E", X"E8E", X"E8D", X"E8D", X"E8C", 
X"E8B", X"E8B", X"E8A", X"E8A", X"E89", X"E89", X"E88", X"E88", 
X"E88", X"E87", X"E87", X"E87", X"E86", X"E86", X"E86", X"E86", 
X"E86", X"E85", X"E85", X"E85", X"E85", X"E85", X"E85", X"E85", 
X"E85", X"E85", X"E85", X"E85", X"E85", X"E85", X"E85", X"E85", 
X"E86", X"E86", X"E86", X"E86", X"E86", X"E87", X"E87", X"E87", 
X"E88", X"E88", X"E88", X"E89", X"E89", X"E8A", X"E8A", X"E8B", 
X"E8B", X"E8C", X"E8D", X"E8D", X"E8E", X"E8E", X"E8F", X"E90", 
X"E91", X"E91", X"E92", X"E93", X"E94", X"E94", X"E95", X"E96", 
X"E97", X"E98", X"E99", X"E9A", X"E9B", X"E9C", X"E9D", X"E9E", 
X"EA0", X"EA1", X"EA2", X"EA3", X"EA4", X"EA6", X"EA7", X"EA8", 
X"EA9", X"EAB", X"EAC", X"EAE", X"EAF", X"EB1", X"EB2", X"EB4", 
X"EB5", X"EB7", X"EB8", X"EBA", X"EBC", X"EBD", X"EBF", X"EC1", 
X"EC3", X"EC4", X"EC6", X"EC8", X"ECA", X"ECC", X"ECE", X"ED0", 
X"ED2", X"ED4", X"ED6", X"ED8", X"EDA", X"EDD", X"EDF", X"EE1", 
X"EE3", X"EE6", X"EE8", X"EEA", X"EED", X"EEF", X"EF2", X"EF4", 
X"EF7", X"EF9", X"EFC", X"EFE", X"F01", X"F03", X"F06", X"F09", 
X"F0C", X"F0F", X"F11", X"F14", X"F17", X"F1A", X"F1D", X"F20", 
X"F23", X"F26", X"F29", X"F2C", X"F30", X"F33", X"F36", X"F39", 
X"F3D", X"F40", X"F43", X"F47", X"F4A", X"F4E", X"F51", X"F54", 
X"F58", X"F5C", X"F5F", X"F63", X"F67", X"F6A", X"F6E", X"F72", 
X"F76", X"F7A", X"F7E", X"F82", X"F85", X"F89", X"F8D", X"F91", 
X"F95", X"F99", X"F9E", X"FA2", X"FA6", X"FAA", X"FAE", X"FB3", 
X"FB7", X"FBB", X"FC0", X"FC4", X"FC9", X"FCD", X"FD1", X"FD6", 
X"FDB", X"FDF", X"FE4", X"FE8", X"FED", X"FF1", X"FF6", X"FFB", 
X"000", X"005", X"009", X"00E", X"013", X"018", X"01D", X"022", 
X"027", X"02C", X"031", X"036", X"03B", X"040", X"045", X"04A", 
X"04F", X"055", X"05A", X"05F", X"064", X"069", X"06F", X"074", 
X"079", X"07F", X"084", X"089", X"08E", X"094", X"099", X"09F", 
X"0A4", X"0AA", X"0AF", X"0B5", X"0BA", X"0C0", X"0C5", X"0CB", 
X"0D0", X"0D6", X"0DB", X"0E1", X"0E7", X"0EC", X"0F2", X"0F7", 
X"0FD", X"102", X"108", X"10E", X"114", X"119", X"11F", X"124", 
X"12A", X"12F", X"135", X"13B", X"141", X"147", X"14C", X"152", 
X"158", X"15D", X"163", X"168", X"16E", X"174", X"179", X"17F", 
X"185", X"18B", X"190", X"196", X"19C", X"1A1", X"1A7", X"1AC", 
X"1B2", X"1B8", X"1BE", X"1C3", X"1C8", X"1CE", X"1D4", X"1D9", 
X"1DF", X"1E4", X"1EA", X"1F0", X"1F5", X"1FA", X"200", X"206", 
X"20B", X"210", X"216", X"21B", X"220", X"226", X"22B", X"231", 
X"236", X"23B", X"241", X"246", X"24B", X"250", X"256", X"25B", 
X"260", X"265", X"26A", X"270", X"275", X"27A", X"27F", X"284", 
X"289", X"28E", X"293", X"298", X"29D", X"2A2", X"2A6", X"2AB", 
X"2B0", X"2B5", X"2BA", X"2BE", X"2C3", X"2C8", X"2CD", X"2D1", 
X"2D6", X"2DA", X"2DF", X"2E3", X"2E8", X"2EC", X"2F1", X"2F5", 
X"2FA", X"2FE", X"302", X"306", X"30B", X"30F", X"313", X"318", 
X"31C", X"320", X"324", X"328", X"32C", X"330", X"334", X"338", 
X"33C", X"340", X"344", X"347", X"34B", X"34F", X"353", X"356", 
X"35A", X"35E", X"361", X"365", X"368", X"36C", X"36F", X"373", 
X"376", X"379", X"37D", X"380", X"384", X"387", X"38A", X"38D", 
X"390", X"394", X"397", X"39A", X"39D", X"3A0", X"3A3", X"3A6", 
X"3A9", X"3AC", X"3AF", X"3B1", X"3B4", X"3B7", X"3BA", X"3BC", 
X"3BF", X"3C2", X"3C4", X"3C7", X"3C9", X"3CC", X"3CF", X"3D1", 
X"3D3", X"3D6", X"3D8", X"3DB", X"3DD", X"3DF", X"3E2", X"3E4", 
X"3E6", X"3E9", X"3EB", X"3ED", X"3EF", X"3F1", X"3F3", X"3F6", 
X"3F8", X"3FA", X"3FC", X"3FE", X"400", X"401", X"403", X"405", 
X"407", X"409", X"40B", X"40D", X"40F", X"410", X"412", X"414", 
X"416", X"417", X"419", X"41B", X"41C", X"41E", X"41F", X"421", 
X"423", X"424", X"426", X"427", X"429", X"42A", X"42C", X"42D", 
X"42F", X"430", X"431", X"433", X"434", X"436", X"437", X"438", 
X"43A", X"43B", X"43C", X"43D", X"43F", X"440", X"441", X"443", 
X"444", X"445", X"446", X"447", X"448", X"44A", X"44B", X"44C", 
X"44D", X"44E", X"44F", X"451", X"452", X"453", X"454", X"455", 
X"456", X"457", X"458", X"459", X"45A", X"45B", X"45C", X"45D", 
X"45F", X"460", X"461", X"462", X"463", X"464", X"465", X"466", 
X"467", X"468", X"469", X"46A", X"46B", X"46C", X"46C", X"46D", 
X"46E", X"46F", X"470", X"471", X"472", X"473", X"474", X"475", 
X"476", X"477", X"478", X"479", X"47A", X"47B", X"47C", X"47D", 
X"47E", X"47F", X"480", X"481", X"481", X"482", X"483", X"484", 
X"485", X"486", X"487", X"488", X"489", X"48A", X"48B", X"48C", 
X"48D", X"48E", X"48F", X"490", X"490", X"491", X"492", X"493", 
X"494", X"495", X"496", X"497", X"498", X"499", X"49A", X"49B", 
X"49C", X"49D", X"49E", X"49F", X"4A0", X"4A1", X"4A2", X"4A2", 
X"4A3", X"4A4", X"4A5", X"4A6", X"4A7", X"4A8", X"4A9", X"4AA", 
X"4AB", X"4AC", X"4AD", X"4AE", X"4AF", X"4B0", X"4B1", X"4B2", 
X"4B3", X"4B4", X"4B5", X"4B6", X"4B7", X"4B8", X"4B9", X"4BA", 
X"4BB", X"4BC", X"4BD", X"4BE", X"4BF", X"4C0", X"4C1", X"4C2", 
X"4C3", X"4C4", X"4C5", X"4C6", X"4C7", X"4C8", X"4C9", X"4CA", 
X"4CB", X"4CC", X"4CD", X"4CE", X"4CF", X"4D0", X"4D1", X"4D2", 
X"4D3", X"4D4", X"4D5", X"4D6", X"4D7", X"4D8", X"4D9", X"4DA", 
X"4DB", X"4DC", X"4DD", X"4DE", X"4DF", X"4E0", X"4E1", X"4E2", 
X"4E3", X"4E4", X"4E5", X"4E6", X"4E7", X"4E9", X"4EA", X"4EB", 
X"4EC", X"4ED", X"4EE", X"4EF", X"4F0", X"4F1", X"4F2", X"4F3", 
X"4F4", X"4F5", X"4F6", X"4F7", X"4F8", X"4F9", X"4FA", X"4FC", 
X"4FD", X"4FE", X"4FF", X"500", X"501", X"502", X"503", X"504", 
X"505", X"506", X"507", X"509", X"50A", X"50B", X"50C", X"50D", 
X"50E", X"50F", X"510", X"512", X"513", X"514", X"515", X"516", 
X"517", X"518", X"519", X"51B", X"51C", X"51D", X"51E", X"51F", 
X"520", X"522", X"523", X"524", X"525", X"526", X"528", X"529", 
X"52A", X"52B", X"52C", X"52E", X"52F", X"530", X"531", X"533", 
X"534", X"535", X"536", X"538", X"539", X"53A", X"53B", X"53D", 
X"53E", X"53F", X"541", X"542", X"543", X"544", X"546", X"547", 
X"548", X"54A", X"54B", X"54C", X"54E", X"54F", X"550", X"552", 
X"553", X"554", X"556", X"557", X"559", X"55A", X"55B", X"55D", 
X"55E", X"55F", X"561", X"562", X"564", X"565", X"567", X"568", 
X"569", X"56B", X"56C", X"56E", X"56F", X"571", X"572", X"573", 
X"575", X"576", X"578", X"579", X"57B", X"57C", X"57E", X"57F", 
X"580", X"582", X"583", X"585", X"586", X"588", X"589", X"58A", 
X"58C", X"58D", X"58F", X"590", X"592", X"593", X"595", X"596", 
X"597", X"599", X"59A", X"59C", X"59D", X"59E", X"5A0", X"5A1", 
X"5A2", X"5A4", X"5A5", X"5A7", X"5A8", X"5A9", X"5AB", X"5AC", 
X"5AD", X"5AE", X"5B0", X"5B1", X"5B2", X"5B3", X"5B5", X"5B6", 
X"5B7", X"5B8", X"5BA", X"5BB", X"5BC", X"5BD", X"5BE", X"5BF", 
X"5C0", X"5C1", X"5C2", X"5C3", X"5C4", X"5C5", X"5C6", X"5C7", 
X"5C8", X"5C9", X"5CA", X"5CB", X"5CC", X"5CC", X"5CD", X"5CE", 
X"5CF", X"5CF", X"5D0", X"5D1", X"5D1", X"5D2", X"5D2", X"5D3", 
X"5D3", X"5D4", X"5D4", X"5D5", X"5D5", X"5D5", X"5D6", X"5D6", 
X"5D6", X"5D6", X"5D6", X"5D6", X"5D6", X"5D6", X"5D6", X"5D6", 
X"5D6", X"5D6", X"5D6", X"5D5", X"5D5", X"5D5", X"5D4", X"5D4", 
X"5D4", X"5D3", X"5D2", X"5D2", X"5D1", X"5D0", X"5D0", X"5CF", 
X"5CE", X"5CD", X"5CC", X"5CB", X"5CA", X"5C9", X"5C7", X"5C6", 
X"5C5", X"5C3", X"5C2", X"5C0", X"5BF", X"5BD", X"5BB", X"5BA", 
X"5B8", X"5B6", X"5B4", X"5B2", X"5B0", X"5AE", X"5AB", X"5A9", 
X"5A7", X"5A4", X"5A2", X"59F", X"59D", X"59A", X"597", X"594", 
X"591", X"58E", X"58B", X"588", X"585", X"582", X"57E", X"57B", 
X"577", X"574", X"570", X"56C", X"568", X"565", X"561", X"55C", 
X"558", X"554", X"550", X"54B", X"547", X"543", X"53E", X"539", 
X"534", X"52F", X"52B", X"525", X"520", X"51B", X"516", X"511", 
X"50B", X"505", X"500", X"4FA", X"4F4", X"4EE", X"4E9", X"4E3", 
X"4DC", X"4D6", X"4D0", X"4CA", X"4C3", X"4BC", X"4B6", X"4AF", 
X"4A8", X"4A1", X"49A", X"494", X"48C", X"485", X"47E", X"476", 
X"46F", X"467", X"460", X"458", X"450", X"448", X"440", X"438", 
X"430", X"428", X"420", X"417", X"40F", X"406", X"3FE", X"3F5", 
X"3EC", X"3E3", X"3DA", X"3D1", X"3C8", X"3BF", X"3B6", X"3AC", 
X"3A3", X"39A", X"390", X"386", X"37C", X"372", X"369", X"35F", 
X"355", X"34B", X"341", X"337", X"32C", X"322", X"318", X"30D", 
X"303", X"2F8", X"2EE", X"2E3", X"2D8", X"2CD", X"2C2", X"2B7", 
X"2AC", X"2A1", X"295", X"28B", X"27F", X"274", X"268", X"25E", 
X"252", X"246", X"23A", X"22E", X"224", X"218", X"20B", X"1FF", 
X"1F4", X"1E8", X"1DC", X"1D0", X"1C4", X"1B8", X"1AC", X"19F", 
X"194", X"187", X"17B", X"16E", X"162", X"156", X"149", X"13D", 
X"130", X"124", X"118", X"10B", X"0FE", X"0F2", X"0E5", X"0D8", 
X"0CC", X"0BF", X"0B3", X"0A6", X"099", X"08C", X"080", X"073", 
X"066", X"059", X"04D", X"040", X"033", X"026", X"01A", X"00D", 
X"000", X"FF2", X"FE5", X"FD9", X"FCC", X"FBF", X"FB2", X"FA6", 
X"F99", X"F8C", X"F7F", X"F73", X"F66", X"F59", X"F4C", X"F40", 
X"F33", X"F27", X"F1A", X"F0D", X"F01", X"EF4", X"EE7", X"EDB", 
X"ECF", X"EC2", X"EB6", X"EA9", X"E9D", X"E91", X"E84", X"E78", 
X"E6B", X"E60", X"E53", X"E47", X"E3B", X"E2F", X"E23", X"E17", 
X"E0B", X"E00", X"DF4", X"DE7", X"DDB", X"DD1", X"DC5", X"DB9", 
X"DAD", X"DA1", X"D97", X"D8B", X"D80", X"D74", X"D6A", X"D5E", 
X"D53", X"D48", X"D3D", X"D32", X"D27", X"D1C", X"D11", X"D07", 
X"CFC", X"CF2", X"CE7", X"CDD", X"CD3", X"CC8", X"CBE", X"CB4", 
X"CAA", X"CA0", X"C96", X"C8D", X"C83", X"C79", X"C6F", X"C65", 
X"C5C", X"C53", X"C49", X"C40", X"C37", X"C2E", X"C25", X"C1C", 
X"C13", X"C0A", X"C01", X"BF9", X"BF0", X"BE8", X"BDF", X"BD7", 
X"BCF", X"BC7", X"BBF", X"BB7", X"BAF", X"BA7", X"B9F", X"B98", 
X"B90", X"B89", X"B81", X"B7A", X"B73", X"B6B", X"B65", X"B5E", 
X"B57", X"B50", X"B49", X"B43", X"B3C", X"B35", X"B2F", X"B29", 
X"B23", X"B1C", X"B16", X"B11", X"B0B", X"B05", X"AFF", X"AFA", 
X"AF4", X"AEE", X"AE9", X"AE4", X"ADF", X"ADA", X"AD4", X"AD0", 
X"ACB", X"AC6", X"AC1", X"ABC", X"AB8", X"AB4", X"AAF", X"AAB", 
X"AA7", X"AA3", X"A9E", X"A9A", X"A97", X"A93", X"A8F", X"A8B", 
X"A88", X"A84", X"A81", X"A7D", X"A7A", X"A77", X"A74", X"A71", 
X"A6E", X"A6B", X"A68", X"A65", X"A62", X"A60", X"A5D", X"A5B", 
X"A58", X"A56", X"A54", X"A51", X"A4F", X"A4D", X"A4B", X"A49", 
X"A47", X"A45", X"A44", X"A42", X"A40", X"A3F", X"A3D", X"A3C", 
X"A3A", X"A39", X"A38", X"A36", X"A35", X"A34", X"A33", X"A32", 
X"A31", X"A30", X"A2F", X"A2F", X"A2E", X"A2D", X"A2D", X"A2C", 
X"A2B", X"A2B", X"A2B", X"A2A", X"A2A", X"A2A", X"A29", X"A29", 
X"A29", X"A29", X"A29", X"A29", X"A29", X"A29", X"A29", X"A29", 
X"A29", X"A29", X"A29", X"A2A", X"A2A", X"A2A", X"A2B", X"A2B", 
X"A2C", X"A2C", X"A2D", X"A2D", X"A2E", X"A2E", X"A2F", X"A30", 
X"A30", X"A31", X"A32", X"A33", X"A33", X"A34", X"A35", X"A36", 
X"A37", X"A38", X"A39", X"A3A", X"A3B", X"A3C", X"A3D", X"A3E", 
X"A3F", X"A40", X"A41", X"A42", X"A43", X"A44", X"A45", X"A47", 
X"A48", X"A49", X"A4A", X"A4C", X"A4D", X"A4E", X"A4F", X"A51", 
X"A52", X"A53", X"A54", X"A56", X"A57", X"A58", X"A5A", X"A5B", 
X"A5D", X"A5E", X"A5F", X"A61", X"A62", X"A63", X"A65", X"A66", 
X"A68", X"A69", X"A6A", X"A6C", X"A6D", X"A6F", X"A70", X"A72", 
X"A73", X"A75", X"A76", X"A77", X"A79", X"A7A", X"A7C", X"A7D", 
X"A7F", X"A80", X"A81", X"A83", X"A84", X"A86", X"A87", X"A89", 
X"A8A", X"A8C", X"A8D", X"A8E", X"A90", X"A91", X"A93", X"A94", 
X"A96", X"A97", X"A98", X"A9A", X"A9B", X"A9D", X"A9E", X"AA0", 
X"AA1", X"AA2", X"AA4", X"AA5", X"AA6", X"AA8", X"AA9", X"AAB", 
X"AAC", X"AAD", X"AAF", X"AB0", X"AB1", X"AB3", X"AB4", X"AB5", 
X"AB7", X"AB8", X"AB9", X"ABB", X"ABC", X"ABD", X"ABE", X"AC0", 
X"AC1", X"AC2", X"AC4", X"AC5", X"AC6", X"AC7", X"AC9", X"ACA", 
X"ACB", X"ACC", X"ACE", X"ACF", X"AD0", X"AD1", X"AD3", X"AD4", 
X"AD5", X"AD6", X"AD7", X"AD9", X"ADA", X"ADB", X"ADC", X"ADD", 
X"ADF", X"AE0", X"AE1", X"AE2", X"AE3", X"AE4", X"AE6", X"AE7", 
X"AE8", X"AE9", X"AEA", X"AEB", X"AEC", X"AED", X"AEF", X"AF0", 
X"AF1", X"AF2", X"AF3", X"AF4", X"AF5", X"AF6", X"AF8", X"AF9", 
X"AFA", X"AFB", X"AFC", X"AFD", X"AFE", X"AFF", X"B00", X"B01", 
X"B02", X"B03", X"B05", X"B06", X"B07", X"B08", X"B09", X"B0A", 
X"B0B", X"B0C", X"B0D", X"B0E", X"B0F", X"B10", X"B11", X"B12", 
X"B13", X"B14", X"B15", X"B16", X"B18", X"B19", X"B1A", X"B1B", 
X"B1C", X"B1D", X"B1E", X"B1F", X"B20", X"B21", X"B22", X"B23", 
X"B24", X"B25", X"B26", X"B27", X"B28", X"B29", X"B2A", X"B2B", 
X"B2C", X"B2D", X"B2E", X"B2F", X"B30", X"B31", X"B32", X"B33", 
X"B34", X"B35", X"B36", X"B37", X"B38", X"B39", X"B3A", X"B3B", 
X"B3C", X"B3D", X"B3E", X"B3F", X"B40", X"B41", X"B42", X"B43", 
X"B44", X"B45", X"B46", X"B47", X"B48", X"B49", X"B4A", X"B4B", 
X"B4C", X"B4D", X"B4E", X"B4F", X"B50", X"B51", X"B52", X"B53", 
X"B54", X"B55", X"B56", X"B57", X"B58", X"B59", X"B5A", X"B5B", 
X"B5C", X"B5D", X"B5D", X"B5E", X"B5F", X"B60", X"B61", X"B62", 
X"B63", X"B64", X"B65", X"B66", X"B67", X"B68", X"B69", X"B6A", 
X"B6B", X"B6C", X"B6D", X"B6E", X"B6F", X"B6F", X"B70", X"B71", 
X"B72", X"B73", X"B74", X"B75", X"B76", X"B77", X"B78", X"B79", 
X"B7A", X"B7B", X"B7C", X"B7D", X"B7E", X"B7E", X"B7F", X"B80", 
X"B81", X"B82", X"B83", X"B84", X"B85", X"B86", X"B87", X"B88", 
X"B89", X"B8A", X"B8B", X"B8C", X"B8D", X"B8E", X"B8F", X"B90", 
X"B91", X"B92", X"B93", X"B93", X"B94", X"B95", X"B96", X"B97", 
X"B98", X"B99", X"B9A", X"B9B", X"B9C", X"B9D", X"B9E", X"B9F", 
X"BA0", X"BA2", X"BA3", X"BA4", X"BA5", X"BA6", X"BA7", X"BA8", 
X"BA9", X"BAA", X"BAB", X"BAC", X"BAD", X"BAE", X"BB0", X"BB1", 
X"BB2", X"BB3", X"BB4", X"BB5", X"BB7", X"BB8", X"BB9", X"BBA", 
X"BBB", X"BBC", X"BBE", X"BBF", X"BC0", X"BC2", X"BC3", X"BC4", 
X"BC5", X"BC7", X"BC8", X"BC9", X"BCB", X"BCC", X"BCE", X"BCF", 
X"BD0", X"BD2", X"BD3", X"BD5", X"BD6", X"BD8", X"BD9", X"BDB", 
X"BDC", X"BDE", X"BE0", X"BE1", X"BE3", X"BE4", X"BE6", X"BE8", 
X"BE9", X"BEB", X"BED", X"BEF", X"BF0", X"BF2", X"BF4", X"BF6", 
X"BF8", X"BFA", X"BFC", X"BFE", X"BFF", X"C01", X"C03", X"C05", 
X"C07", X"C09", X"C0C", X"C0E", X"C10", X"C12", X"C14", X"C16", 
X"C19", X"C1B", X"C1D", X"C20", X"C22", X"C24", X"C27", X"C29", 
X"C2C", X"C2E", X"C30", X"C33", X"C36", X"C38", X"C3B", X"C3D", 
X"C40", X"C43", X"C45", X"C48", X"C4B", X"C4E", X"C50", X"C53", 
X"C56", X"C59", X"C5C", X"C5F", X"C62", X"C65", X"C68", X"C6B", 
X"C6F", X"C72", X"C75", X"C78", X"C7B", X"C7F", X"C82", X"C86", 
X"C89", X"C8C", X"C90", X"C93", X"C97", X"C9A", X"C9E", X"CA1", 
X"CA5", X"CA9", X"CAC", X"CB0", X"CB4", X"CB8", X"CBB", X"CBF", 
X"CC3", X"CC7", X"CCB", X"CCF", X"CD3", X"CD7", X"CDB", X"CDF", 
X"CE3", X"CE7", X"CEC", X"CF0", X"CF4", X"CF9", X"CFD", X"D01", 
X"D05", X"D0A", X"D0E", X"D13", X"D17", X"D1C", X"D20", X"D25", 
X"D29", X"D2E", X"D32", X"D37", X"D3C", X"D41", X"D45", X"D4A", 
X"D4F", X"D54", X"D59", X"D5D", X"D62", X"D67", X"D6C", X"D71", 
X"D76", X"D7B", X"D80", X"D85", X"D8A", X"D8F", X"D95", X"D9A", 
X"D9F", X"DA4", X"DA9", X"DAF", X"DB4", X"DB9", X"DBE", X"DC4", 
X"DC9", X"DCE", X"DD4", X"DD9", X"DDF", X"DE4", X"DE9", X"DEF", 
X"DF4", X"DF9", X"DFF", X"E05", X"E0A", X"E0F", X"E15", X"E1B", 
X"E20", X"E26", X"E2B", X"E31", X"E37", X"E3C", X"E41", X"E47", 
X"E4D", X"E53", X"E58", X"E5E", X"E63", X"E69", X"E6F", X"E74", 
X"E7A", X"E80", X"E86", X"E8B", X"E91", X"E97", X"E9C", X"EA2", 
X"EA7", X"EAD", X"EB3", X"EB8", X"EBE", X"EC4", X"ECA", X"ED0", 
X"ED5", X"EDB", X"EE0", X"EE6", X"EEB", X"EF1", X"EF7", X"EFD", 
X"F02", X"F08", X"F0D", X"F13", X"F18", X"F1E", X"F24", X"F29", 
X"F2F", X"F34", X"F3A", X"F3F", X"F45", X"F4A", X"F50", X"F55", 
X"F5B", X"F60", X"F66", X"F6B", X"F71", X"F76", X"F7B", X"F80", 
X"F86", X"F8B", X"F90", X"F96", X"F9B", X"FA0", X"FA5", X"FAA", 
X"FB0", X"FB5", X"FBA", X"FBF", X"FC4", X"FC9", X"FCE", X"FD3", 
X"FD8", X"FDD", X"FE2", X"FE7", X"FEC", X"FF1", X"FF6", X"FFA", 
X"FFF", X"004", X"009", X"00E", X"012", X"017", X"01B", X"020", 
X"024", X"029", X"02E", X"032", X"036", X"03B", X"03F", X"044", 
X"048", X"04C", X"051", X"055", X"059", X"05D", X"061", X"066", 
X"06A", X"06E", X"072", X"076", X"07A", X"07D", X"081", X"085", 
X"089", X"08D", X"091", X"095", X"098", X"09C", X"0A0", X"0A3", 
X"0A7", X"0AB", X"0AE", X"0B1", X"0B5", X"0B8", X"0BC", X"0BF", 
X"0C2", X"0C6", X"0C9", X"0CC", X"0CF", X"0D3", X"0D6", X"0D9", 
X"0DC", X"0DF", X"0E2", X"0E5", X"0E8", X"0EB", X"0EE", X"0F0", 
X"0F3", X"0F6", X"0F9", X"0FC", X"0FE", X"101", X"103", X"106", 
X"108", X"10B", X"10D", X"110", X"112", X"115", X"117", X"119", 
X"11C", X"11E", X"120", X"122", X"125", X"127", X"129", X"12B", 
X"12D", X"12F", X"131", X"133", X"135", X"137", X"139", X"13B", 
X"13C", X"13E", X"140", X"142", X"143", X"145", X"147", X"148", 
X"14A", X"14B", X"14D", X"14E", X"150", X"151", X"153", X"154", 
X"156", X"157", X"158", X"159", X"15B", X"15C", X"15D", X"15E", 
X"15F", X"161", X"162", X"163", X"164", X"165", X"166", X"167", 
X"168", X"169", X"16A", X"16B", X"16B", X"16C", X"16D", X"16E", 
X"16E", X"16F", X"170", X"171", X"171", X"172", X"172", X"173", 
X"174", X"174", X"175", X"175", X"176", X"176", X"177", X"177", 
X"177", X"178", X"178", X"178", X"179", X"179", X"179", X"179", 
X"179", X"17A", X"17A", X"17A", X"17A", X"17A", X"17A", X"17A", 
X"17A", X"17A", X"17A", X"17A", X"17A", X"17A", X"17A", X"17A", 
X"179", X"179", X"179", X"179", X"179", X"178", X"178", X"178", 
X"177", X"177", X"177", X"176", X"176", X"175", X"175", X"174", 
X"174", X"173", X"172", X"172", X"171", X"171", X"170", X"16F", 
X"16E", X"16E", X"16D", X"16C", X"16B", X"16B", X"16A", X"169", 
X"168", X"167", X"166", X"165", X"164", X"163", X"162", X"161", 
X"15F", X"15E", X"15D", X"15C", X"15B", X"159", X"158", X"157", 
X"156", X"154", X"153", X"151", X"150", X"14E", X"14D", X"14B", 
X"14A", X"148", X"147", X"145", X"143", X"142", X"140", X"13E", 
X"13C", X"13B", X"139", X"137", X"135", X"133", X"131", X"12F", 
X"12D", X"12B", X"129", X"127", X"125", X"122", X"120", X"11E", 
X"11C", X"119", X"117", X"115", X"112", X"110", X"10D", X"10B", 
X"108", X"106", X"103", X"101", X"0FE", X"0FC", X"0F9", X"0F6", 
X"0F3", X"0F0", X"0EE", X"0EB", X"0E8", X"0E5", X"0E2", X"0DF", 
X"0DC", X"0D9", X"0D6", X"0D3", X"0CF", X"0CC", X"0C9", X"0C6", 
X"0C2", X"0BF", X"0BC", X"0B8", X"0B5", X"0B1", X"0AE", X"0AB", 
X"0A7", X"0A3", X"0A0", X"09C", X"098", X"095", X"091", X"08D", 
X"089", X"085", X"081", X"07D", X"07A", X"076", X"072", X"06E", 
X"06A", X"066", X"061", X"05D", X"059", X"055", X"051", X"04C", 
X"048", X"044", X"03F", X"03B", X"036", X"032", X"02E", X"029", 
X"024", X"020", X"01B", X"017", X"012", X"00E", X"009", X"004", 
X"FFF", X"FFA", X"FF6", X"FF1", X"FEC", X"FE7", X"FE2", X"FDD", 
X"FD8", X"FD3", X"FCE", X"FC9", X"FC4", X"FBF", X"FBA", X"FB5", 
X"FB0", X"FAA", X"FA5", X"FA0", X"F9B", X"F96", X"F90", X"F8B", 
X"F86", X"F80", X"F7B", X"F76", X"F71", X"F6B", X"F66", X"F60", 
X"F5B", X"F55", X"F50", X"F4A", X"F45", X"F3F", X"F3A", X"F34", 
X"F2F", X"F29", X"F24", X"F1E", X"F18", X"F13", X"F0D", X"F08", 
X"F02", X"EFD", X"EF7", X"EF1", X"EEB", X"EE6", X"EE0", X"EDB", 
X"ED5", X"ED0", X"ECA", X"EC4", X"EBE", X"EB8", X"EB3", X"EAD", 
X"EA7", X"EA2", X"E9C", X"E97", X"E91", X"E8B", X"E86", X"E80", 
X"E7A", X"E74", X"E6F", X"E69", X"E63", X"E5E", X"E58", X"E53", 
X"E4D", X"E47", X"E41", X"E3C", X"E37", X"E31", X"E2B", X"E26", 
X"E20", X"E1B", X"E15", X"E0F", X"E0A", X"E05", X"DFF", X"DF9", 
X"DF4", X"DEF", X"DE9", X"DE4", X"DDF", X"DD9", X"DD4", X"DCE", 
X"DC9", X"DC4", X"DBE", X"DB9", X"DB4", X"DAF", X"DA9", X"DA4", 
X"D9F", X"D9A", X"D95", X"D8F", X"D8A", X"D85", X"D80", X"D7B", 
X"D76", X"D71", X"D6C", X"D67", X"D62", X"D5D", X"D59", X"D54", 
X"D4F", X"D4A", X"D45", X"D41", X"D3C", X"D37", X"D32", X"D2E", 
X"D29", X"D25", X"D20", X"D1C", X"D17", X"D13", X"D0E", X"D0A", 
X"D05", X"D01", X"CFD", X"CF9", X"CF4", X"CF0", X"CEC", X"CE7", 
X"CE3", X"CDF", X"CDB", X"CD7", X"CD3", X"CCF", X"CCB", X"CC7", 
X"CC3", X"CBF", X"CBB", X"CB8", X"CB4", X"CB0", X"CAC", X"CA9", 
X"CA5", X"CA1", X"C9E", X"C9A", X"C97", X"C93", X"C90", X"C8C", 
X"C89", X"C86", X"C82", X"C7F", X"C7B", X"C78", X"C75", X"C72", 
X"C6F", X"C6B", X"C68", X"C65", X"C62", X"C5F", X"C5C", X"C59", 
X"C56", X"C53", X"C50", X"C4E", X"C4B", X"C48", X"C45", X"C43", 
X"C40", X"C3D", X"C3B", X"C38", X"C36", X"C33", X"C30", X"C2E", 
X"C2C", X"C29", X"C27", X"C24", X"C22", X"C20", X"C1D", X"C1B", 
X"C19", X"C16", X"C14", X"C12", X"C10", X"C0E", X"C0C", X"C09", 
X"C07", X"C05", X"C03", X"C01", X"BFF", X"BFE", X"BFC", X"BFA", 
X"BF8", X"BF6", X"BF4", X"BF2", X"BF0", X"BEF", X"BED", X"BEB", 
X"BE9", X"BE8", X"BE6", X"BE4", X"BE3", X"BE1", X"BE0", X"BDE", 
X"BDC", X"BDB", X"BD9", X"BD8", X"BD6", X"BD5", X"BD3", X"BD2", 
X"BD0", X"BCF", X"BCE", X"BCC", X"BCB", X"BC9", X"BC8", X"BC7", 
X"BC5", X"BC4", X"BC3", X"BC2", X"BC0", X"BBF", X"BBE", X"BBC", 
X"BBB", X"BBA", X"BB9", X"BB8", X"BB7", X"BB5", X"BB4", X"BB3", 
X"BB2", X"BB1", X"BB0", X"BAE", X"BAD", X"BAC", X"BAB", X"BAA", 
X"BA9", X"BA8", X"BA7", X"BA6", X"BA5", X"BA4", X"BA3", X"BA2", 
X"BA0", X"B9F", X"B9E", X"B9D", X"B9C", X"B9B", X"B9A", X"B99", 
X"B98", X"B97", X"B96", X"B95", X"B94", X"B93", X"B93", X"B92", 
X"B91", X"B90", X"B8F", X"B8E", X"B8D", X"B8C", X"B8B", X"B8A", 
X"B89", X"B88", X"B87", X"B86", X"B85", X"B84", X"B83", X"B82", 
X"B81", X"B80", X"B7F", X"B7E", X"B7E", X"B7D", X"B7C", X"B7B", 
X"B7A", X"B79", X"B78", X"B77", X"B76", X"B75", X"B74", X"B73", 
X"B72", X"B71", X"B70", X"B6F", X"B6F", X"B6E", X"B6D", X"B6C", 
X"B6B", X"B6A", X"B69", X"B68", X"B67", X"B66", X"B65", X"B64", 
X"B63", X"B62", X"B61", X"B60", X"B5F", X"B5E", X"B5D", X"B5D", 
X"B5C", X"B5B", X"B5A", X"B59", X"B58", X"B57", X"B56", X"B55", 
X"B54", X"B53", X"B52", X"B51", X"B50", X"B4F", X"B4E", X"B4D", 
X"B4C", X"B4B", X"B4A", X"B49", X"B48", X"B47", X"B46", X"B45", 
X"B44", X"B43", X"B42", X"B41", X"B40", X"B3F", X"B3E", X"B3D", 
X"B3C", X"B3B", X"B3A", X"B39", X"B38", X"B37", X"B36", X"B35", 
X"B34", X"B33", X"B32", X"B31", X"B30", X"B2F", X"B2E", X"B2D", 
X"B2C", X"B2B", X"B2A", X"B29", X"B28", X"B27", X"B26", X"B25", 
X"B24", X"B23", X"B22", X"B21", X"B20", X"B1F", X"B1E", X"B1D", 
X"B1C", X"B1B", X"B1A", X"B19", X"B18", X"B16", X"B15", X"B14", 
X"B13", X"B12", X"B11", X"B10", X"B0F", X"B0E", X"B0D", X"B0C", 
X"B0B", X"B0A", X"B09", X"B08", X"B07", X"B06", X"B05", X"B03", 
X"B02", X"B01", X"B00", X"AFF", X"AFE", X"AFD", X"AFC", X"AFB", 
X"AFA", X"AF9", X"AF8", X"AF6", X"AF5", X"AF4", X"AF3", X"AF2", 
X"AF1", X"AF0", X"AEF", X"AED", X"AEC", X"AEB", X"AEA", X"AE9", 
X"AE8", X"AE7", X"AE6", X"AE4", X"AE3", X"AE2", X"AE1", X"AE0", 
X"ADF", X"ADD", X"ADC", X"ADB", X"ADA", X"AD9", X"AD7", X"AD6", 
X"AD5", X"AD4", X"AD3", X"AD1", X"AD0", X"ACF", X"ACE", X"ACC", 
X"ACB", X"ACA", X"AC9", X"AC7", X"AC6", X"AC5", X"AC4", X"AC2", 
X"AC1", X"AC0", X"ABE", X"ABD", X"ABC", X"ABB", X"AB9", X"AB8", 
X"AB7", X"AB5", X"AB4", X"AB3", X"AB1", X"AB0", X"AAF", X"AAD", 
X"AAC", X"AAB", X"AA9", X"AA8", X"AA6", X"AA5", X"AA4", X"AA2", 
X"AA1", X"AA0", X"A9E", X"A9D", X"A9B", X"A9A", X"A98", X"A97", 
X"A96", X"A94", X"A93", X"A91", X"A90", X"A8E", X"A8D", X"A8C", 
X"A8A", X"A89", X"A87", X"A86", X"A84", X"A83", X"A81", X"A80", 
X"A7F", X"A7D", X"A7C", X"A7A", X"A79", X"A77", X"A76", X"A75", 
X"A73", X"A72", X"A70", X"A6F", X"A6D", X"A6C", X"A6A", X"A69", 
X"A68", X"A66", X"A65", X"A63", X"A62", X"A61", X"A5F", X"A5E", 
X"A5D", X"A5B", X"A5A", X"A58", X"A57", X"A56", X"A54", X"A53", 
X"A52", X"A51", X"A4F", X"A4E", X"A4D", X"A4C", X"A4A", X"A49", 
X"A48", X"A47", X"A45", X"A44", X"A43", X"A42", X"A41", X"A40", 
X"A3F", X"A3E", X"A3D", X"A3C", X"A3B", X"A3A", X"A39", X"A38", 
X"A37", X"A36", X"A35", X"A34", X"A33", X"A33", X"A32", X"A31", 
X"A30", X"A30", X"A2F", X"A2E", X"A2E", X"A2D", X"A2D", X"A2C", 
X"A2C", X"A2B", X"A2B", X"A2A", X"A2A", X"A2A", X"A29", X"A29", 
X"A29", X"A29", X"A29", X"A29", X"A29", X"A29", X"A29", X"A29", 
X"A29", X"A29", X"A29", X"A2A", X"A2A", X"A2A", X"A2B", X"A2B", 
X"A2B", X"A2C", X"A2D", X"A2D", X"A2E", X"A2F", X"A2F", X"A30", 
X"A31", X"A32", X"A33", X"A34", X"A35", X"A36", X"A38", X"A39", 
X"A3A", X"A3C", X"A3D", X"A3F", X"A40", X"A42", X"A44", X"A45", 
X"A47", X"A49", X"A4B", X"A4D", X"A4F", X"A51", X"A54", X"A56", 
X"A58", X"A5B", X"A5D", X"A60", X"A62", X"A65", X"A68", X"A6B", 
X"A6E", X"A71", X"A74", X"A77", X"A7A", X"A7D", X"A81", X"A84", 
X"A88", X"A8B", X"A8F", X"A93", X"A97", X"A9A", X"A9E", X"AA3", 
X"AA7", X"AAB", X"AAF", X"AB4", X"AB8", X"ABC", X"AC1", X"AC6", 
X"ACB", X"AD0", X"AD4", X"ADA", X"ADF", X"AE4", X"AE9", X"AEE", 
X"AF4", X"AFA", X"AFF", X"B05", X"B0B", X"B11", X"B16", X"B1C", 
X"B23", X"B29", X"B2F", X"B35", X"B3C", X"B43", X"B49", X"B50", 
X"B57", X"B5E", X"B65", X"B6B", X"B73", X"B7A", X"B81", X"B89", 
X"B90", X"B98", X"B9F", X"BA7", X"BAF", X"BB7", X"BBF", X"BC7", 
X"BCF", X"BD7", X"BDF", X"BE8", X"BF0", X"BF9", X"C01", X"C0A", 
X"C13", X"C1C", X"C25", X"C2E", X"C37", X"C40", X"C49", X"C53", 
X"C5C", X"C65", X"C6F", X"C79", X"C83", X"C8D", X"C96", X"CA0", 
X"CAA", X"CB4", X"CBE", X"CC8", X"CD3", X"CDD", X"CE7", X"CF2", 
X"CFC", X"D07", X"D11", X"D1C", X"D27", X"D32", X"D3D", X"D48", 
X"D53", X"D5E", X"D6A", X"D74", X"D80", X"D8B", X"D97", X"DA1", 
X"DAD", X"DB9", X"DC5", X"DD1", X"DDB", X"DE7", X"DF4", X"E00", 
X"E0B", X"E17", X"E23", X"E2F", X"E3B", X"E47", X"E53", X"E60", 
X"E6B", X"E78", X"E84", X"E91", X"E9D", X"EA9", X"EB6", X"EC2", 
X"ECF", X"EDB", X"EE7", X"EF4", X"F01", X"F0D", X"F1A", X"F27", 
X"F33", X"F40", X"F4C", X"F59", X"F66", X"F73", X"F7F", X"F8C", 
X"F99", X"FA6", X"FB2", X"FBF", X"FCC", X"FD9", X"FE5", X"FF2" 
);

signal data : std_logic_vector(31 downto 0);
signal unsignedIndex : unsigned(11 downto 0) := X"000";

begin

rom_select: process (clk, en)
begin
	if (rising_edge(clk)) then
    if (en = '1') then
		unsignedIndex <= unsigned(address_reg);
		data <= (SIN_ROM(to_integer(unsignedIndex)) & x"00000");
		sin_out <= std_logic_vector(shift_right(signed(data), 20));
    end if;
  end if;
end process rom_select;

end rtl;
