  --------------------------------------------------------------------------------------------------------------------------
-- Original Authors : Simon Doherty, Eric Lunty, Kyle Brooks, Peter Roland						--
-- Date created: N/A 													--
--															--
-- Additional Authors : Randi Derbyshire, Adam Narten, Oliver Rarog, Celeste Chiasson					--
-- Date edited: March 26, 2018											--
--															--
-- This program takes a value from the synthesizer.vhd file and runs it through the 12-bit ROM to find the 	 	--
-- respective sine wave value. 												--
--------------------------------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use IEEE.STD_LOGIC_SIGNED.all;
use ieee.numeric_std.all;               -- Needed for shifts

entity HarpSin_lut is

port (
	clk      : in  std_logic;
	en       : in  std_logic;
	
	--Address input
	address_reg : in std_logic_vector(11 downto 0); 
	
	--Sine value output
	sin_out  : out std_logic_vector(31 downto 0)
	);
end entity;


architecture rtl of HarpSin_lut is


type rom_type is array (0 to 4095) of std_logic_vector (11 downto 0);

constant SIN_ROM : rom_type :=

(
X"000", X"00D", X"01A", X"026", X"033", X"040", X"04D", X"059", 
X"066", X"073", X"080", X"08C", X"099", X"0A6", X"0B3", X"0BE", 
X"0CB", X"0D8", X"0E5", X"0F2", X"0FE", X"10B", X"117", X"124", 
X"130", X"13D", X"149", X"156", X"162", X"16E", X"17B", X"187", 
X"194", X"19F", X"1AC", X"1B8", X"1C4", X"1D0", X"1DC", X"1E8", 
X"1F4", X"1FF", X"20B", X"218", X"224", X"22E", X"23A", X"246", 
X"252", X"25E", X"269", X"274", X"280", X"28B", X"296", X"2A1", 
X"2AD", X"2B8", X"2C2", X"2CD", X"2D9", X"2E4", X"2EF", X"2F9", 
X"303", X"30E", X"319", X"323", X"32D", X"338", X"342", X"34C", 
X"356", X"361", X"36B", X"374", X"37E", X"388", X"392", X"39C", 
X"3A5", X"3AF", X"3B8", X"3C2", X"3CA", X"3D4", X"3DD", X"3E6", 
X"3EF", X"3F8", X"401", X"40A", X"413", X"41B", X"423", X"42C", 
X"434", X"43C", X"445", X"44D", X"455", X"45C", X"465", X"46D", 
X"474", X"47C", X"483", X"48B", X"493", X"49A", X"4A1", X"4A8", 
X"4AF", X"4B7", X"4BD", X"4C4", X"4CB", X"4D2", X"4D8", X"4DF", 
X"4E5", X"4EC", X"4F2", X"4F8", X"4FE", X"504", X"50A", X"510", 
X"516", X"51C", X"521", X"527", X"52C", X"532", X"537", X"53C", 
X"542", X"547", X"54C", X"551", X"556", X"55B", X"55F", X"564", 
X"568", X"56D", X"572", X"576", X"57A", X"57E", X"583", X"587", 
X"58B", X"58F", X"593", X"597", X"59B", X"59E", X"5A2", X"5A5", 
X"5A9", X"5AC", X"5B0", X"5B3", X"5B6", X"5B9", X"5BC", X"5C0", 
X"5C3", X"5C6", X"5C8", X"5CB", X"5CE", X"5D1", X"5D3", X"5D6", 
X"5D9", X"5DB", X"5DD", X"5E0", X"5E2", X"5E5", X"5E7", X"5E9", 
X"5EB", X"5ED", X"5EF", X"5F1", X"5F3", X"5F5", X"5F7", X"5F9", 
X"5FB", X"5FD", X"5FE", X"600", X"602", X"603", X"605", X"606", 
X"608", X"609", X"60B", X"60C", X"60D", X"60F", X"610", X"611", 
X"612", X"614", X"615", X"616", X"617", X"618", X"619", X"61A", 
X"61C", X"61C", X"61D", X"61E", X"61F", X"620", X"621", X"622", 
X"623", X"624", X"625", X"626", X"626", X"627", X"628", X"629", 
X"62A", X"62A", X"62B", X"62C", X"62D", X"62D", X"62E", X"62F", 
X"630", X"630", X"631", X"632", X"632", X"633", X"634", X"635", 
X"635", X"636", X"637", X"638", X"638", X"639", X"63A", X"63A", 
X"63B", X"63C", X"63D", X"63E", X"63E", X"63F", X"640", X"641", 
X"641", X"642", X"643", X"644", X"645", X"646", X"647", X"647", 
X"648", X"649", X"64A", X"64B", X"64C", X"64D", X"64E", X"64F", 
X"650", X"651", X"652", X"653", X"654", X"655", X"657", X"658", 
X"659", X"65A", X"65B", X"65C", X"65E", X"65F", X"660", X"661", 
X"663", X"664", X"665", X"667", X"668", X"66A", X"66B", X"66C", 
X"66E", X"66F", X"671", X"672", X"674", X"676", X"677", X"679", 
X"67A", X"67C", X"67E", X"67F", X"681", X"683", X"684", X"686", 
X"688", X"68A", X"68B", X"68D", X"68F", X"691", X"693", X"695", 
X"697", X"699", X"69A", X"69C", X"69F", X"6A0", X"6A2", X"6A4", 
X"6A7", X"6A8", X"6AA", X"6AD", X"6AF", X"6B1", X"6B3", X"6B5", 
X"6B7", X"6B9", X"6BB", X"6BE", X"6C0", X"6C2", X"6C4", X"6C6", 
X"6C8", X"6CB", X"6CD", X"6CF", X"6D1", X"6D4", X"6D6", X"6D8", 
X"6DA", X"6DC", X"6DF", X"6E1", X"6E3", X"6E5", X"6E8", X"6EA", 
X"6EC", X"6EE", X"6F1", X"6F3", X"6F5", X"6F7", X"6FA", X"6FC", 
X"6FE", X"700", X"703", X"705", X"707", X"709", X"70B", X"70D", 
X"70F", X"712", X"714", X"716", X"718", X"71A", X"71C", X"71E", 
X"720", X"722", X"724", X"726", X"728", X"72A", X"72C", X"72E", 
X"730", X"732", X"734", X"736", X"738", X"739", X"73B", X"73D", 
X"73F", X"740", X"742", X"744", X"745", X"747", X"748", X"74A", 
X"74B", X"74D", X"74E", X"750", X"751", X"753", X"754", X"755", 
X"756", X"758", X"759", X"75A", X"75B", X"75C", X"75D", X"75E", 
X"75F", X"760", X"761", X"762", X"763", X"763", X"764", X"765", 
X"765", X"766", X"767", X"767", X"768", X"768", X"768", X"769", 
X"769", X"769", X"76A", X"76A", X"76A", X"76A", X"76A", X"76A", 
X"76A", X"76A", X"76A", X"769", X"769", X"769", X"769", X"768", 
X"768", X"767", X"767", X"766", X"765", X"765", X"764", X"763", 
X"762", X"761", X"761", X"760", X"75F", X"75D", X"75C", X"75B", 
X"75A", X"759", X"757", X"756", X"755", X"753", X"751", X"750", 
X"74E", X"74D", X"74B", X"749", X"747", X"745", X"743", X"742", 
X"740", X"73D", X"73B", X"739", X"737", X"735", X"732", X"730", 
X"72E", X"72B", X"729", X"726", X"724", X"721", X"71E", X"71B", 
X"718", X"716", X"713", X"710", X"70D", X"70A", X"707", X"704", 
X"701", X"6FE", X"6FB", X"6F7", X"6F4", X"6F1", X"6ED", X"6EA", 
X"6E6", X"6E3", X"6E0", X"6DC", X"6D8", X"6D5", X"6D1", X"6CD", 
X"6CA", X"6C6", X"6C2", X"6BE", X"6BA", X"6B6", X"6B3", X"6AF", 
X"6AB", X"6A6", X"6A2", X"69F", X"69A", X"696", X"692", X"68E", 
X"68A", X"685", X"681", X"67D", X"679", X"674", X"670", X"66B", 
X"667", X"663", X"65E", X"65A", X"656", X"651", X"64C", X"648", 
X"644", X"63F", X"63A", X"636", X"632", X"62D", X"628", X"623", 
X"61F", X"61A", X"616", X"611", X"60C", X"608", X"603", X"5FE", 
X"5FA", X"5F5", X"5F1", X"5EC", X"5E7", X"5E2", X"5DE", X"5D9", 
X"5D4", X"5D0", X"5CB", X"5C7", X"5C2", X"5BD", X"5B9", X"5B4", 
X"5AF", X"5AB", X"5A6", X"5A2", X"59D", X"598", X"594", X"58F", 
X"58B", X"586", X"581", X"57D", X"579", X"574", X"570", X"56B", 
X"567", X"562", X"55E", X"559", X"555", X"551", X"54D", X"548", 
X"544", X"540", X"53C", X"537", X"534", X"52F", X"52B", X"527", 
X"523", X"51F", X"51B", X"517", X"513", X"50F", X"50B", X"507", 
X"503", X"500", X"4FC", X"4F8", X"4F4", X"4F1", X"4ED", X"4E9", 
X"4E6", X"4E2", X"4DF", X"4DB", X"4D8", X"4D4", X"4D1", X"4CE", 
X"4CA", X"4C7", X"4C4", X"4C1", X"4BD", X"4BA", X"4B7", X"4B4", 
X"4B1", X"4AE", X"4AB", X"4A8", X"4A5", X"4A3", X"4A0", X"49D", 
X"49A", X"498", X"495", X"493", X"490", X"48D", X"48B", X"488", 
X"486", X"484", X"481", X"47F", X"47D", X"47B", X"478", X"476", 
X"474", X"472", X"470", X"46E", X"46C", X"46A", X"469", X"467", 
X"465", X"463", X"462", X"460", X"45E", X"45D", X"45B", X"45A", 
X"458", X"457", X"455", X"454", X"453", X"451", X"450", X"44F", 
X"44E", X"44D", X"44C", X"44B", X"44A", X"449", X"448", X"447", 
X"446", X"445", X"444", X"443", X"443", X"442", X"441", X"441", 
X"440", X"43F", X"43F", X"43E", X"43E", X"43D", X"43D", X"43C", 
X"43C", X"43C", X"43B", X"43B", X"43B", X"43B", X"43A", X"43A", 
X"43A", X"43A", X"43A", X"43A", X"43A", X"439", X"439", X"439", 
X"439", X"43A", X"43A", X"43A", X"43A", X"43A", X"43A", X"43A", 
X"43A", X"43B", X"43B", X"43B", X"43B", X"43B", X"43C", X"43C", 
X"43C", X"43D", X"43D", X"43D", X"43E", X"43E", X"43E", X"43F", 
X"43F", X"440", X"440", X"440", X"441", X"441", X"442", X"442", 
X"443", X"443", X"444", X"444", X"445", X"445", X"445", X"446", 
X"446", X"447", X"447", X"448", X"448", X"449", X"449", X"44A", 
X"44A", X"44B", X"44B", X"44C", X"44C", X"44D", X"44D", X"44E", 
X"44E", X"44E", X"44F", X"44F", X"450", X"450", X"451", X"451", 
X"451", X"452", X"452", X"453", X"453", X"453", X"454", X"454", 
X"454", X"454", X"455", X"455", X"455", X"456", X"456", X"456", 
X"456", X"456", X"457", X"457", X"457", X"457", X"457", X"457", 
X"457", X"457", X"457", X"457", X"457", X"457", X"457", X"457", 
X"457", X"457", X"457", X"457", X"457", X"456", X"456", X"456", 
X"456", X"456", X"455", X"455", X"455", X"454", X"454", X"454", 
X"453", X"453", X"452", X"452", X"451", X"451", X"450", X"450", 
X"44F", X"44F", X"44E", X"44D", X"44D", X"44C", X"44B", X"44B", 
X"44A", X"449", X"448", X"447", X"447", X"446", X"445", X"444", 
X"443", X"442", X"441", X"440", X"43F", X"43E", X"43D", X"43C", 
X"43B", X"439", X"438", X"437", X"436", X"435", X"434", X"432", 
X"431", X"430", X"42E", X"42D", X"42C", X"42A", X"429", X"427", 
X"426", X"424", X"423", X"421", X"420", X"41E", X"41D", X"41B", 
X"41A", X"418", X"416", X"415", X"413", X"411", X"40F", X"40E", 
X"40C", X"40A", X"408", X"407", X"405", X"403", X"401", X"3FF", 
X"3FD", X"3FC", X"3FA", X"3F8", X"3F6", X"3F4", X"3F2", X"3F0", 
X"3EE", X"3EC", X"3EA", X"3E8", X"3E6", X"3E3", X"3E2", X"3DF", 
X"3DD", X"3DB", X"3D9", X"3D7", X"3D5", X"3D2", X"3D0", X"3CE", 
X"3CC", X"3CA", X"3C8", X"3C5", X"3C3", X"3C1", X"3BF", X"3BC", 
X"3BA", X"3B8", X"3B5", X"3B3", X"3B1", X"3AF", X"3AC", X"3AA", 
X"3A8", X"3A5", X"3A3", X"3A0", X"39E", X"39C", X"399", X"397", 
X"395", X"392", X"390", X"38D", X"38B", X"389", X"386", X"384", 
X"382", X"37F", X"37D", X"37A", X"378", X"375", X"373", X"370", 
X"36E", X"36C", X"369", X"367", X"364", X"362", X"35F", X"35D", 
X"35A", X"358", X"355", X"353", X"350", X"34E", X"34B", X"349", 
X"346", X"344", X"341", X"33F", X"33C", X"33A", X"337", X"335", 
X"332", X"330", X"32D", X"32B", X"328", X"326", X"323", X"321", 
X"31E", X"31C", X"319", X"317", X"314", X"311", X"30F", X"30D", 
X"30A", X"307", X"305", X"302", X"300", X"2FD", X"2FA", X"2F8", 
X"2F5", X"2F3", X"2F0", X"2EE", X"2EB", X"2E9", X"2E6", X"2E3", 
X"2E1", X"2DE", X"2DC", X"2D9", X"2D6", X"2D4", X"2D1", X"2CE", 
X"2CC", X"2C9", X"2C7", X"2C4", X"2C1", X"2BF", X"2BC", X"2B9", 
X"2B7", X"2B4", X"2B1", X"2AF", X"2AC", X"2A9", X"2A6", X"2A4", 
X"2A1", X"29E", X"29C", X"299", X"296", X"293", X"290", X"28E", 
X"28B", X"288", X"285", X"282", X"27F", X"27C", X"27A", X"277", 
X"274", X"271", X"26E", X"26B", X"268", X"265", X"262", X"25F", 
X"25C", X"259", X"256", X"253", X"250", X"24D", X"24A", X"247", 
X"244", X"241", X"23E", X"23A", X"237", X"234", X"231", X"22E", 
X"22A", X"227", X"224", X"221", X"21D", X"21A", X"217", X"213", 
X"210", X"20D", X"209", X"206", X"202", X"1FF", X"1FC", X"1F8", 
X"1F4", X"1F1", X"1EE", X"1EA", X"1E6", X"1E3", X"1DF", X"1DB", 
X"1D8", X"1D4", X"1D0", X"1CD", X"1C9", X"1C5", X"1C1", X"1BE", 
X"1BA", X"1B6", X"1B2", X"1AE", X"1AA", X"1A6", X"1A2", X"19E", 
X"19A", X"196", X"192", X"18E", X"18A", X"186", X"182", X"17D", 
X"17A", X"175", X"171", X"16D", X"169", X"164", X"160", X"15C", 
X"157", X"153", X"14F", X"14A", X"146", X"141", X"13D", X"138", 
X"134", X"130", X"12B", X"126", X"122", X"11D", X"119", X"114", 
X"10F", X"10A", X"106", X"101", X"0FC", X"0F7", X"0F3", X"0EE", 
X"0E9", X"0E4", X"0E0", X"0DB", X"0D6", X"0D1", X"0CC", X"0C7", 
X"0C2", X"0BD", X"0B8", X"0B4", X"0AE", X"0A9", X"0A4", X"0A0", 
X"09A", X"095", X"090", X"08B", X"086", X"081", X"07C", X"077", 
X"072", X"06D", X"067", X"062", X"05D", X"058", X"053", X"04D", 
X"049", X"043", X"03E", X"039", X"033", X"02E", X"029", X"024", 
X"01E", X"01A", X"014", X"00F", X"009", X"005", X"FFF", X"FFA", 
X"FF5", X"FF0", X"FEA", X"FE5", X"FE0", X"FDA", X"FD5", X"FD0", 
X"FCB", X"FC5", X"FC1", X"FBB", X"FB6", X"FB1", X"FAC", X"FA7", 
X"FA1", X"F9C", X"F97", X"F92", X"F8D", X"F88", X"F83", X"F7E", 
X"F79", X"F73", X"F6E", X"F6A", X"F65", X"F5F", X"F5A", X"F56", 
X"F51", X"F4C", X"F47", X"F42", X"F3D", X"F38", X"F33", X"F2E", 
X"F2A", X"F25", X"F20", X"F1C", X"F17", X"F12", X"F0E", X"F09", 
X"F04", X"F00", X"EFB", X"EF7", X"EF2", X"EEE", X"EEA", X"EE5", 
X"EE1", X"EDD", X"ED8", X"ED4", X"ED0", X"ECC", X"EC8", X"EC3", 
X"EBF", X"EBB", X"EB7", X"EB3", X"EAF", X"EAB", X"EA8", X"EA4", 
X"EA0", X"E9C", X"E99", X"E95", X"E91", X"E8D", X"E8A", X"E86", 
X"E83", X"E7F", X"E7C", X"E79", X"E75", X"E72", X"E6F", X"E6C", 
X"E69", X"E65", X"E62", X"E60", X"E5D", X"E5A", X"E57", X"E54", 
X"E51", X"E4E", X"E4C", X"E49", X"E46", X"E44", X"E41", X"E3F", 
X"E3D", X"E3A", X"E38", X"E35", X"E33", X"E31", X"E2F", X"E2D", 
X"E2B", X"E29", X"E27", X"E25", X"E23", X"E22", X"E20", X"E1E", 
X"E1C", X"E1B", X"E19", X"E18", X"E16", X"E15", X"E14", X"E12", 
X"E11", X"E10", X"E0F", X"E0E", X"E0D", X"E0C", X"E0B", X"E0A", 
X"E09", X"E08", X"E07", X"E07", X"E06", X"E05", X"E05", X"E04", 
X"E04", X"E03", X"E03", X"E03", X"E02", X"E02", X"E02", X"E02", 
X"E02", X"E01", X"E01", X"E02", X"E02", X"E02", X"E02", X"E02", 
X"E02", X"E03", X"E03", X"E03", X"E04", X"E04", X"E05", X"E05", 
X"E06", X"E06", X"E07", X"E08", X"E08", X"E09", X"E0A", X"E0B", 
X"E0C", X"E0C", X"E0D", X"E0E", X"E0F", X"E10", X"E11", X"E13", 
X"E14", X"E15", X"E16", X"E17", X"E19", X"E1A", X"E1B", X"E1D", 
X"E1E", X"E1F", X"E21", X"E22", X"E24", X"E25", X"E27", X"E28", 
X"E2A", X"E2B", X"E2D", X"E2F", X"E30", X"E32", X"E34", X"E35", 
X"E37", X"E39", X"E3B", X"E3C", X"E3E", X"E40", X"E42", X"E44", 
X"E46", X"E48", X"E49", X"E4B", X"E4D", X"E4F", X"E51", X"E53", 
X"E55", X"E57", X"E59", X"E5B", X"E5D", X"E5F", X"E61", X"E63", 
X"E65", X"E67", X"E69", X"E6B", X"E6D", X"E6F", X"E71", X"E73", 
X"E75", X"E77", X"E79", X"E7B", X"E7D", X"E7F", X"E81", X"E83", 
X"E85", X"E87", X"E88", X"E8A", X"E8C", X"E8E", X"E90", X"E92", 
X"E94", X"E96", X"E98", X"E99", X"E9B", X"E9D", X"E9F", X"EA1", 
X"EA2", X"EA4", X"EA6", X"EA8", X"EA9", X"EAB", X"EAD", X"EAE", 
X"EB0", X"EB2", X"EB3", X"EB5", X"EB7", X"EB8", X"EBA", X"EBB", 
X"EBD", X"EBE", X"EC0", X"EC1", X"EC2", X"EC4", X"EC5", X"EC6", 
X"EC8", X"EC9", X"ECA", X"ECC", X"ECD", X"ECE", X"ECF", X"ED0", 
X"ED1", X"ED2", X"ED3", X"ED4", X"ED5", X"ED6", X"ED7", X"ED8", 
X"ED9", X"EDA", X"EDB", X"EDC", X"EDC", X"EDD", X"EDE", X"EDE", 
X"EDF", X"EE0", X"EE0", X"EE1", X"EE1", X"EE2", X"EE2", X"EE3", 
X"EE3", X"EE4", X"EE4", X"EE5", X"EE5", X"EE5", X"EE5", X"EE6", 
X"EE6", X"EE6", X"EE6", X"EE6", X"EE6", X"EE6", X"EE7", X"EE7", 
X"EE7", X"EE7", X"EE6", X"EE6", X"EE6", X"EE6", X"EE6", X"EE6", 
X"EE6", X"EE5", X"EE5", X"EE5", X"EE5", X"EE4", X"EE4", X"EE3", 
X"EE3", X"EE3", X"EE2", X"EE2", X"EE1", X"EE1", X"EE0", X"EE0", 
X"EDF", X"EDF", X"EDE", X"EDE", X"EDD", X"EDC", X"EDC", X"EDB", 
X"EDA", X"EDA", X"ED9", X"ED8", X"ED7", X"ED7", X"ED6", X"ED5", 
X"ED4", X"ED4", X"ED3", X"ED2", X"ED1", X"ED0", X"ECF", X"ECF", 
X"ECE", X"ECD", X"ECC", X"ECB", X"ECA", X"EC9", X"EC9", X"EC8", 
X"EC7", X"EC6", X"EC5", X"EC4", X"EC3", X"EC2", X"EC2", X"EC1", 
X"EC0", X"EBF", X"EBE", X"EBD", X"EBD", X"EBC", X"EBB", X"EBA", 
X"EB9", X"EB8", X"EB8", X"EB7", X"EB6", X"EB5", X"EB4", X"EB4", 
X"EB3", X"EB2", X"EB2", X"EB1", X"EB0", X"EB0", X"EAF", X"EAE", 
X"EAE", X"EAD", X"EAD", X"EAC", X"EAC", X"EAB", X"EAB", X"EAA", 
X"EAA", X"EA9", X"EA9", X"EA9", X"EA8", X"EA8", X"EA8", X"EA8", 
X"EA7", X"EA7", X"EA7", X"EA7", X"EA7", X"EA7", X"EA7", X"EA7", 
X"EA7", X"EA7", X"EA7", X"EA7", X"EA7", X"EA7", X"EA8", X"EA8", 
X"EA8", X"EA8", X"EA9", X"EA9", X"EAA", X"EAA", X"EAB", X"EAB", 
X"EAC", X"EAC", X"EAD", X"EAE", X"EAF", X"EAF", X"EB0", X"EB1", 
X"EB2", X"EB3", X"EB4", X"EB5", X"EB6", X"EB7", X"EB8", X"EBA", 
X"EBB", X"EBC", X"EBD", X"EBF", X"EC0", X"EC2", X"EC3", X"EC5", 
X"EC6", X"EC8", X"ECA", X"ECC", X"ECD", X"ECF", X"ED1", X"ED3", 
X"ED5", X"ED7", X"ED9", X"EDB", X"EDD", X"EDF", X"EE2", X"EE4", 
X"EE6", X"EE9", X"EEB", X"EED", X"EF0", X"EF2", X"EF5", X"EF8", 
X"EFA", X"EFD", X"F00", X"F03", X"F05", X"F08", X"F0B", X"F0E", 
X"F11", X"F14", X"F17", X"F1A", X"F1D", X"F21", X"F24", X"F27", 
X"F2A", X"F2E", X"F31", X"F35", X"F38", X"F3B", X"F3F", X"F43", 
X"F46", X"F4A", X"F4E", X"F51", X"F55", X"F59", X"F5C", X"F60", 
X"F64", X"F68", X"F6C", X"F70", X"F74", X"F78", X"F7C", X"F80", 
X"F84", X"F88", X"F8C", X"F90", X"F95", X"F99", X"F9D", X"FA1", 
X"FA5", X"FAA", X"FAE", X"FB2", X"FB7", X"FBB", X"FC0", X"FC4", 
X"FC8", X"FCD", X"FD1", X"FD5", X"FDA", X"FDE", X"FE3", X"FE7", 
X"FEB", X"FF0", X"FF5", X"FF9", X"FFD", X"002", X"006", X"00B", 
X"00F", X"014", X"018", X"01D", X"021", X"026", X"02A", X"02F", 
X"033", X"038", X"03C", X"041", X"045", X"049", X"04E", X"052", 
X"057", X"05B", X"05F", X"064", X"068", X"06D", X"071", X"075", 
X"079", X"07E", X"081", X"086", X"08A", X"08E", X"092", X"096", 
X"09A", X"09E", X"0A2", X"0A6", X"0AA", X"0AE", X"0B2", X"0B6", 
X"0B9", X"0BD", X"0C1", X"0C5", X"0C8", X"0CC", X"0D0", X"0D3", 
X"0D7", X"0DA", X"0DE", X"0E1", X"0E4", X"0E7", X"0EB", X"0EE", 
X"0F1", X"0F4", X"0F7", X"0FA", X"0FD", X"100", X"103", X"106", 
X"108", X"10B", X"10E", X"110", X"113", X"115", X"118", X"11A", 
X"11D", X"11F", X"121", X"123", X"125", X"127", X"129", X"12B", 
X"12D", X"12F", X"130", X"132", X"134", X"135", X"137", X"138", 
X"13A", X"13B", X"13C", X"13D", X"13E", X"13F", X"140", X"141", 
X"142", X"143", X"143", X"144", X"145", X"145", X"146", X"146", 
X"146", X"146", X"147", X"147", X"147", X"147", X"147", X"146", 
X"146", X"146", X"145", X"145", X"144", X"144", X"143", X"142", 
X"142", X"141", X"140", X"13F", X"13E", X"13D", X"13C", X"13A", 
X"139", X"138", X"136", X"135", X"133", X"131", X"130", X"12E", 
X"12C", X"12A", X"128", X"126", X"124", X"122", X"120", X"11D", 
X"11B", X"119", X"116", X"114", X"111", X"10E", X"10C", X"109", 
X"106", X"103", X"101", X"0FE", X"0FA", X"0F7", X"0F4", X"0F1", 
X"0EE", X"0EA", X"0E7", X"0E4", X"0E0", X"0DD", X"0D9", X"0D6", 
X"0D2", X"0CF", X"0CB", X"0C7", X"0C3", X"0BF", X"0BB", X"0B7", 
X"0B4", X"0B0", X"0AC", X"0A7", X"0A4", X"09F", X"09B", X"097", 
X"093", X"08F", X"08A", X"086", X"081", X"07D", X"079", X"074", 
X"070", X"06B", X"067", X"062", X"05D", X"059", X"055", X"050", 
X"04B", X"046", X"042", X"03D", X"038", X"034", X"02F", X"02A", 
X"026", X"021", X"01C", X"017", X"013", X"00E", X"009", X"004", 
X"000", X"FFB", X"FF6", X"FF1", X"FEC", X"FE8", X"FE3", X"FDE", 
X"FD9", X"FD5", X"FD0", X"FCB", X"FC7", X"FC2", X"FBD", X"FB9", 
X"FB4", X"FAF", X"FAA", X"FA6", X"FA2", X"F9D", X"F98", X"F94", 
X"F8F", X"F8B", X"F86", X"F82", X"F7E", X"F79", X"F75", X"F70", 
X"F6C", X"F68", X"F64", X"F60", X"F5B", X"F58", X"F53", X"F4F", 
X"F4B", X"F48", X"F44", X"F40", X"F3C", X"F38", X"F34", X"F30", 
X"F2D", X"F29", X"F26", X"F22", X"F1F", X"F1B", X"F18", X"F15", 
X"F11", X"F0E", X"F0B", X"F08", X"F05", X"F01", X"EFE", X"EFC", 
X"EF9", X"EF6", X"EF3", X"EF1", X"EEE", X"EEB", X"EE9", X"EE6", 
X"EE4", X"EE2", X"EDF", X"EDD", X"EDB", X"ED9", X"ED7", X"ED5", 
X"ED3", X"ED1", X"ECF", X"ECE", X"ECC", X"ECA", X"EC9", X"EC7", 
X"EC6", X"EC5", X"EC3", X"EC2", X"EC1", X"EC0", X"EBF", X"EBE", 
X"EBD", X"EBD", X"EBC", X"EBB", X"EBB", X"EBA", X"EBA", X"EB9", 
X"EB9", X"EB9", X"EB8", X"EB8", X"EB8", X"EB8", X"EB8", X"EB9", 
X"EB9", X"EB9", X"EB9", X"EBA", X"EBA", X"EBB", X"EBC", X"EBC", 
X"EBD", X"EBE", X"EBF", X"EC0", X"EC1", X"EC2", X"EC3", X"EC4", 
X"EC5", X"EC7", X"EC8", X"ECA", X"ECB", X"ECD", X"ECF", X"ED0", 
X"ED2", X"ED4", X"ED6", X"ED8", X"EDA", X"EDC", X"EDE", X"EE0", 
X"EE2", X"EE5", X"EE7", X"EEA", X"EEC", X"EEF", X"EF1", X"EF4", 
X"EF7", X"EF9", X"EFC", X"EFF", X"F02", X"F05", X"F08", X"F0B", 
X"F0E", X"F11", X"F14", X"F18", X"F1B", X"F1E", X"F21", X"F25", 
X"F28", X"F2C", X"F2F", X"F33", X"F37", X"F3A", X"F3E", X"F42", 
X"F46", X"F49", X"F4D", X"F51", X"F55", X"F59", X"F5D", X"F61", 
X"F65", X"F69", X"F6D", X"F71", X"F75", X"F79", X"F7E", X"F81", 
X"F86", X"F8A", X"F8E", X"F92", X"F97", X"F9B", X"FA0", X"FA4", 
X"FA8", X"FAD", X"FB1", X"FB6", X"FBA", X"FBE", X"FC3", X"FC7", 
X"FCC", X"FD0", X"FD5", X"FD9", X"FDE", X"FE2", X"FE7", X"FEB", 
X"FF0", X"FF4", X"FF9", X"FFD", X"002", X"006", X"00A", X"00F", 
X"014", X"018", X"01C", X"021", X"025", X"02A", X"02E", X"032", 
X"037", X"03B", X"03F", X"044", X"048", X"04D", X"051", X"055", 
X"05A", X"05E", X"062", X"066", X"06A", X"06F", X"073", X"077", 
X"07B", X"07F", X"083", X"087", X"08B", X"08F", X"093", X"097", 
X"09B", X"09F", X"0A3", X"0A6", X"0AA", X"0AE", X"0B1", X"0B5", 
X"0B9", X"0BC", X"0C0", X"0C4", X"0C7", X"0CA", X"0CE", X"0D1", 
X"0D5", X"0D8", X"0DB", X"0DE", X"0E2", X"0E5", X"0E8", X"0EB", 
X"0EE", X"0F1", X"0F4", X"0F7", X"0FA", X"0FC", X"0FF", X"102", 
X"105", X"107", X"10A", X"10D", X"10F", X"112", X"114", X"116", 
X"119", X"11B", X"11D", X"120", X"122", X"124", X"126", X"128", 
X"12A", X"12C", X"12E", X"130", X"132", X"133", X"135", X"137", 
X"139", X"13A", X"13C", X"13D", X"13F", X"140", X"142", X"143", 
X"144", X"145", X"147", X"148", X"149", X"14A", X"14B", X"14C", 
X"14D", X"14E", X"14F", X"150", X"150", X"151", X"152", X"153", 
X"153", X"154", X"154", X"155", X"155", X"156", X"156", X"157", 
X"157", X"157", X"157", X"158", X"158", X"158", X"158", X"158", 
X"158", X"158", X"158", X"158", X"158", X"158", X"158", X"158", 
X"158", X"157", X"157", X"157", X"157", X"156", X"156", X"156", 
X"155", X"155", X"154", X"154", X"153", X"153", X"152", X"152", 
X"151", X"151", X"150", X"14F", X"14F", X"14E", X"14D", X"14D", 
X"14C", X"14B", X"14B", X"14A", X"149", X"148", X"147", X"147", 
X"146", X"145", X"144", X"143", X"142", X"142", X"141", X"140", 
X"13F", X"13E", X"13D", X"13D", X"13C", X"13B", X"13A", X"139", 
X"138", X"137", X"136", X"136", X"135", X"134", X"133", X"132", 
X"131", X"130", X"130", X"12F", X"12E", X"12D", X"12C", X"12B", 
X"12B", X"12A", X"129", X"128", X"128", X"127", X"126", X"125", 
X"125", X"124", X"123", X"123", X"122", X"121", X"121", X"120", 
X"120", X"11F", X"11F", X"11E", X"11E", X"11D", X"11D", X"11C", 
X"11C", X"11C", X"11B", X"11B", X"11A", X"11A", X"11A", X"11A", 
X"119", X"119", X"119", X"119", X"119", X"119", X"119", X"118", 
X"118", X"118", X"118", X"119", X"119", X"119", X"119", X"119", 
X"119", X"119", X"11A", X"11A", X"11A", X"11A", X"11B", X"11B", 
X"11C", X"11C", X"11D", X"11D", X"11E", X"11E", X"11F", X"11F", 
X"120", X"121", X"121", X"122", X"123", X"123", X"124", X"125", 
X"126", X"127", X"128", X"129", X"12A", X"12B", X"12C", X"12D", 
X"12E", X"12F", X"130", X"131", X"132", X"133", X"135", X"136", 
X"137", X"139", X"13A", X"13B", X"13D", X"13E", X"13F", X"141", 
X"142", X"144", X"145", X"147", X"148", X"14A", X"14C", X"14D", 
X"14F", X"151", X"152", X"154", X"156", X"157", X"159", X"15B", 
X"15D", X"15E", X"160", X"162", X"164", X"166", X"167", X"169", 
X"16B", X"16D", X"16F", X"171", X"173", X"175", X"177", X"178", 
X"17A", X"17C", X"17E", X"180", X"182", X"184", X"186", X"188", 
X"18A", X"18C", X"18E", X"190", X"192", X"194", X"196", X"198", 
X"19A", X"19C", X"19E", X"1A0", X"1A2", X"1A4", X"1A6", X"1A8", 
X"1AA", X"1AC", X"1AE", X"1B0", X"1B2", X"1B4", X"1B6", X"1B7", 
X"1B9", X"1BB", X"1BD", X"1BF", X"1C1", X"1C3", X"1C4", X"1C6", 
X"1C8", X"1CA", X"1CB", X"1CD", X"1CF", X"1D0", X"1D2", X"1D4", 
X"1D5", X"1D7", X"1D8", X"1DA", X"1DB", X"1DD", X"1DE", X"1E0", 
X"1E1", X"1E2", X"1E4", X"1E5", X"1E6", X"1E8", X"1E9", X"1EA", 
X"1EB", X"1EC", X"1EE", X"1EF", X"1F0", X"1F1", X"1F2", X"1F3", 
X"1F3", X"1F4", X"1F5", X"1F6", X"1F7", X"1F7", X"1F8", X"1F9", 
X"1F9", X"1FA", X"1FA", X"1FB", X"1FB", X"1FC", X"1FC", X"1FC", 
X"1FD", X"1FD", X"1FD", X"1FD", X"1FD", X"1FD", X"1FE", X"1FE", 
X"1FD", X"1FD", X"1FD", X"1FD", X"1FD", X"1FC", X"1FC", X"1FC", 
X"1FB", X"1FB", X"1FA", X"1FA", X"1F9", X"1F8", X"1F8", X"1F7", 
X"1F6", X"1F5", X"1F4", X"1F3", X"1F2", X"1F1", X"1F0", X"1EF", 
X"1EE", X"1ED", X"1EB", X"1EA", X"1E9", X"1E7", X"1E6", X"1E4", 
X"1E3", X"1E1", X"1DF", X"1DD", X"1DC", X"1DA", X"1D8", X"1D6", 
X"1D4", X"1D2", X"1D0", X"1CE", X"1CC", X"1CA", X"1C7", X"1C5", 
X"1C2", X"1C0", X"1BE", X"1BB", X"1B9", X"1B6", X"1B3", X"1B1", 
X"1AE", X"1AB", X"1A8", X"1A5", X"1A2", X"19F", X"19D", X"19A", 
X"196", X"193", X"190", X"18D", X"18A", X"186", X"183", X"180", 
X"17C", X"179", X"175", X"172", X"16E", X"16A", X"166", X"163", 
X"15F", X"15B", X"157", X"154", X"150", X"14C", X"148", X"144", 
X"140", X"13C", X"137", X"133", X"12F", X"12B", X"127", X"122", 
X"11E", X"11A", X"115", X"111", X"10D", X"108", X"104", X"0FF", 
X"0FB", X"0F6", X"0F1", X"0ED", X"0E8", X"0E3", X"0DF", X"0DA", 
X"0D5", X"0D1", X"0CC", X"0C7", X"0C2", X"0BD", X"0B8", X"0B3", 
X"0AE", X"0A9", X"0A5", X"0A0", X"09A", X"095", X"091", X"08C", 
X"086", X"081", X"07C", X"077", X"072", X"06D", X"068", X"063", 
X"05E", X"058", X"053", X"04E", X"049", X"044", X"03E", X"03A", 
X"034", X"02F", X"02A", X"025", X"01F", X"01A", X"015", X"00F", 
X"00A", X"005", X"000", X"FFA", X"FF6", X"FF0", X"FEB", X"FE5", 
X"FE1", X"FDB", X"FD6", X"FD1", X"FCC", X"FC6", X"FC1", X"FBC", 
X"FB6", X"FB2", X"FAC", X"FA7", X"FA2", X"F9D", X"F98", X"F92", 
X"F8D", X"F88", X"F83", X"F7E", X"F79", X"F74", X"F6F", X"F6A", 
X"F65", X"F5F", X"F5B", X"F56", X"F51", X"F4B", X"F47", X"F42", 
X"F3D", X"F38", X"F33", X"F2E", X"F29", X"F24", X"F1F", X"F1B", 
X"F16", X"F11", X"F0C", X"F08", X"F03", X"EFE", X"EF9", X"EF5", 
X"EF0", X"EEB", X"EE6", X"EE2", X"EDD", X"ED9", X"ED4", X"ECF", 
X"ECB", X"EC7", X"EC2", X"EBE", X"EB9", X"EB5", X"EB0", X"EAC", 
X"EA8", X"EA3", X"E9F", X"E9B", X"E96", X"E92", X"E8E", X"E8A", 
X"E85", X"E82", X"E7D", X"E79", X"E75", X"E71", X"E6D", X"E69", 
X"E65", X"E61", X"E5D", X"E59", X"E55", X"E51", X"E4D", X"E49", 
X"E45", X"E41", X"E3E", X"E3A", X"E36", X"E32", X"E2F", X"E2B", 
X"E27", X"E24", X"E20", X"E1C", X"E19", X"E15", X"E11", X"E0E", 
X"E0B", X"E07", X"E03", X"E00", X"DFD", X"DF9", X"DF6", X"DF2", 
X"DEF", X"DEC", X"DE8", X"DE5", X"DE2", X"DDE", X"DDB", X"DD8", 
X"DD5", X"DD1", X"DCE", X"DCB", X"DC8", X"DC5", X"DC1", X"DBE", 
X"DBB", X"DB8", X"DB5", X"DB2", X"DAF", X"DAC", X"DA9", X"DA6", 
X"DA3", X"DA0", X"D9D", X"D9A", X"D97", X"D94", X"D91", X"D8E", 
X"D8B", X"D88", X"D85", X"D83", X"D80", X"D7D", X"D7A", X"D77", 
X"D74", X"D71", X"D6F", X"D6C", X"D69", X"D66", X"D63", X"D61", 
X"D5E", X"D5B", X"D59", X"D56", X"D53", X"D50", X"D4E", X"D4B", 
X"D48", X"D46", X"D43", X"D40", X"D3E", X"D3B", X"D38", X"D36", 
X"D33", X"D31", X"D2E", X"D2B", X"D29", X"D26", X"D23", X"D21", 
X"D1E", X"D1C", X"D19", X"D16", X"D14", X"D11", X"D0F", X"D0C", 
X"D0A", X"D07", X"D05", X"D02", X"CFF", X"CFD", X"CFA", X"CF8", 
X"CF5", X"CF2", X"CF0", X"CEE", X"CEB", X"CE8", X"CE6", X"CE3", 
X"CE1", X"CDE", X"CDC", X"CD9", X"CD7", X"CD4", X"CD2", X"CCF", 
X"CCD", X"CCA", X"CC8", X"CC5", X"CC3", X"CC0", X"CBE", X"CBB", 
X"CB9", X"CB6", X"CB4", X"CB1", X"CAF", X"CAC", X"CAA", X"CA7", 
X"CA5", X"CA2", X"CA0", X"C9D", X"C9B", X"C98", X"C96", X"C93", 
X"C91", X"C8F", X"C8C", X"C8A", X"C87", X"C85", X"C82", X"C80", 
X"C7D", X"C7B", X"C79", X"C76", X"C74", X"C72", X"C6F", X"C6D", 
X"C6A", X"C68", X"C66", X"C63", X"C61", X"C5F", X"C5C", X"C5A", 
X"C57", X"C55", X"C53", X"C50", X"C4E", X"C4C", X"C4A", X"C47", 
X"C45", X"C43", X"C40", X"C3E", X"C3C", X"C3A", X"C37", X"C35", 
X"C33", X"C31", X"C2F", X"C2D", X"C2A", X"C28", X"C26", X"C24", 
X"C22", X"C20", X"C1D", X"C1C", X"C19", X"C17", X"C15", X"C13", 
X"C11", X"C0F", X"C0D", X"C0B", X"C09", X"C07", X"C05", X"C03", 
X"C02", X"C00", X"BFE", X"BFC", X"BFA", X"BF8", X"BF7", X"BF5", 
X"BF3", X"BF1", X"BF0", X"BEE", X"BEC", X"BEA", X"BE9", X"BE7", 
X"BE5", X"BE4", X"BE2", X"BE1", X"BDF", X"BDE", X"BDC", X"BDB", 
X"BD9", X"BD8", X"BD6", X"BD5", X"BD3", X"BD2", X"BD1", X"BCF", 
X"BCE", X"BCD", X"BCB", X"BCA", X"BC9", X"BC8", X"BC7", X"BC6", 
X"BC4", X"BC3", X"BC2", X"BC1", X"BC0", X"BBF", X"BBE", X"BBD", 
X"BBC", X"BBB", X"BBA", X"BB9", X"BB8", X"BB8", X"BB7", X"BB6", 
X"BB5", X"BB4", X"BB4", X"BB3", X"BB2", X"BB2", X"BB1", X"BB0", 
X"BB0", X"BAF", X"BAF", X"BAE", X"BAE", X"BAD", X"BAD", X"BAC", 
X"BAC", X"BAB", X"BAB", X"BAB", X"BAA", X"BAA", X"BAA", X"BA9", 
X"BA9", X"BA9", X"BA9", X"BA9", X"BA8", X"BA8", X"BA8", X"BA8", 
X"BA8", X"BA8", X"BA8", X"BA8", X"BA8", X"BA8", X"BA8", X"BA8", 
X"BA8", X"BA8", X"BA8", X"BA8", X"BA8", X"BA8", X"BA8", X"BA9", 
X"BA9", X"BA9", X"BA9", X"BA9", X"BAA", X"BAA", X"BAA", X"BAB", 
X"BAB", X"BAB", X"BAB", X"BAC", X"BAC", X"BAC", X"BAD", X"BAD", 
X"BAE", X"BAE", X"BAE", X"BAF", X"BAF", X"BB0", X"BB0", X"BB1", 
X"BB1", X"BB1", X"BB2", X"BB2", X"BB3", X"BB3", X"BB4", X"BB4", 
X"BB5", X"BB5", X"BB6", X"BB6", X"BB7", X"BB7", X"BB8", X"BB8", 
X"BB9", X"BB9", X"BBA", X"BBA", X"BBA", X"BBB", X"BBB", X"BBC", 
X"BBC", X"BBD", X"BBD", X"BBE", X"BBE", X"BBF", X"BBF", X"BBF", 
X"BC0", X"BC0", X"BC1", X"BC1", X"BC1", X"BC2", X"BC2", X"BC2", 
X"BC3", X"BC3", X"BC3", X"BC4", X"BC4", X"BC4", X"BC4", X"BC4", 
X"BC5", X"BC5", X"BC5", X"BC5", X"BC5", X"BC5", X"BC5", X"BC5", 
X"BC6", X"BC6", X"BC6", X"BC6", X"BC5", X"BC5", X"BC5", X"BC5", 
X"BC5", X"BC5", X"BC5", X"BC4", X"BC4", X"BC4", X"BC4", X"BC3", 
X"BC3", X"BC3", X"BC2", X"BC2", X"BC1", X"BC1", X"BC0", X"BC0", 
X"BBF", X"BBE", X"BBE", X"BBD", X"BBC", X"BBC", X"BBB", X"BBA", 
X"BB9", X"BB8", X"BB7", X"BB6", X"BB5", X"BB4", X"BB3", X"BB2", 
X"BB1", X"BB0", X"BAF", X"BAE", X"BAC", X"BAB", X"BAA", X"BA8", 
X"BA7", X"BA5", X"BA4", X"BA2", X"BA1", X"B9F", X"B9D", X"B9C", 
X"B9A", X"B98", X"B96", X"B95", X"B93", X"B91", X"B8F", X"B8D", 
X"B8B", X"B89", X"B87", X"B84", X"B82", X"B80", X"B7E", X"B7B", 
X"B79", X"B77", X"B74", X"B72", X"B6F", X"B6C", X"B6A", X"B67", 
X"B65", X"B62", X"B5F", X"B5C", X"B5A", X"B57", X"B54", X"B51", 
X"B4E", X"B4B", X"B48", X"B45", X"B42", X"B3E", X"B3B", X"B38", 
X"B35", X"B31", X"B2E", X"B2B", X"B27", X"B24", X"B20", X"B1D", 
X"B19", X"B16", X"B12", X"B0E", X"B0B", X"B07", X"B03", X"AFF", 
X"AFC", X"AF8", X"AF4", X"AF0", X"AEC", X"AE8", X"AE4", X"AE0", 
X"ADC", X"AD8", X"AD4", X"AD0", X"ACB", X"AC8", X"AC3", X"ABF", 
X"ABB", X"AB7", X"AB2", X"AAE", X"AAA", X"AA6", X"AA1", X"A9D", 
X"A98", X"A94", X"A8F", X"A8B", X"A86", X"A82", X"A7E", X"A79", 
X"A74", X"A70", X"A6B", X"A67", X"A62", X"A5D", X"A59", X"A54", 
X"A50", X"A4B", X"A46", X"A42", X"A3D", X"A38", X"A34", X"A2F", 
X"A2B", X"A26", X"A21", X"A1D", X"A18", X"A13", X"A0E", X"A0A", 
X"A05", X"A01", X"9FC", X"9F7", X"9F3", X"9EE", X"9E9", X"9E5", 
X"9E0", X"9DC", X"9D7", X"9D2", X"9CD", X"9C9", X"9C5", X"9C0", 
X"9BB", X"9B7", X"9B3", X"9AE", X"9A9", X"9A5", X"9A1", X"99C", 
X"998", X"994", X"98F", X"98B", X"986", X"982", X"97E", X"97A", 
X"975", X"971", X"96D", X"969", X"965", X"960", X"95D", X"959", 
X"954", X"950", X"94C", X"949", X"945", X"941", X"93D", X"939", 
X"935", X"932", X"92E", X"92A", X"927", X"923", X"91F", X"91C", 
X"919", X"915", X"912", X"90E", X"90B", X"908", X"904", X"901", 
X"8FE", X"8FB", X"8F8", X"8F5", X"8F2", X"8EF", X"8EC", X"8E9", 
X"8E6", X"8E4", X"8E1", X"8DE", X"8DB", X"8D9", X"8D6", X"8D4", 
X"8D1", X"8CF", X"8CD", X"8CA", X"8C8", X"8C6", X"8C4", X"8C2", 
X"8BF", X"8BD", X"8BC", X"8BA", X"8B8", X"8B6", X"8B4", X"8B2", 
X"8B1", X"8AF", X"8AE", X"8AC", X"8AA", X"8A9", X"8A8", X"8A6", 
X"8A5", X"8A4", X"8A3", X"8A2", X"8A0", X"89F", X"89E", X"89E", 
X"89D", X"89C", X"89B", X"89A", X"89A", X"899", X"898", X"898", 
X"897", X"897", X"896", X"896", X"896", X"896", X"895", X"895", 
X"895", X"895", X"895", X"895", X"895", X"895", X"895", X"896", 
X"896", X"896", X"897", X"897", X"897", X"898", X"898", X"899", 
X"89A", X"89A", X"89B", X"89C", X"89C", X"89D", X"89E", X"89F", 
X"8A0", X"8A1", X"8A2", X"8A3", X"8A4", X"8A5", X"8A6", X"8A7", 
X"8A9", X"8AA", X"8AB", X"8AC", X"8AE", X"8AF", X"8B1", X"8B2", 
X"8B4", X"8B5", X"8B7", X"8B8", X"8BA", X"8BB", X"8BD", X"8BF", 
X"8C0", X"8C2", X"8C4", X"8C6", X"8C7", X"8C9", X"8CB", X"8CD", 
X"8CF", X"8D1", X"8D3", X"8D5", X"8D7", X"8D9", X"8DB", X"8DD", 
X"8DF", X"8E1", X"8E3", X"8E5", X"8E7", X"8E9", X"8EB", X"8ED", 
X"8F0", X"8F2", X"8F4", X"8F6", X"8F8", X"8FA", X"8FC", X"8FF", 
X"901", X"903", X"905", X"908", X"90A", X"90C", X"90E", X"911", 
X"913", X"915", X"917", X"91A", X"91C", X"91E", X"920", X"923", 
X"925", X"927", X"929", X"92B", X"92E", X"930", X"932", X"934", 
X"937", X"939", X"93B", X"93D", X"93F", X"941", X"944", X"946", 
X"948", X"94A", X"94C", X"94E", X"950", X"952", X"955", X"957", 
X"958", X"95B", X"95D", X"95F", X"960", X"963", X"965", X"966", 
X"968", X"96A", X"96C", X"96E", X"970", X"972", X"974", X"975", 
X"977", X"979", X"97B", X"97C", X"97E", X"980", X"981", X"983", 
X"985", X"986", X"988", X"989", X"98B", X"98D", X"98E", X"990", 
X"991", X"993", X"994", X"995", X"997", X"998", X"99A", X"99B", 
X"99C", X"99E", X"99F", X"9A0", X"9A1", X"9A3", X"9A4", X"9A5", 
X"9A6", X"9A7", X"9A8", X"9AA", X"9AB", X"9AC", X"9AD", X"9AE", 
X"9AF", X"9B0", X"9B1", X"9B2", X"9B3", X"9B4", X"9B5", X"9B6", 
X"9B7", X"9B8", X"9B8", X"9B9", X"9BA", X"9BB", X"9BC", X"9BD", 
X"9BE", X"9BE", X"9BF", X"9C0", X"9C1", X"9C1", X"9C2", X"9C3", 
X"9C4", X"9C5", X"9C5", X"9C6", X"9C7", X"9C7", X"9C8", X"9C9", 
X"9CA", X"9CA", X"9CB", X"9CC", X"9CD", X"9CD", X"9CE", X"9CF", 
X"9CF", X"9D0", X"9D1", X"9D2", X"9D2", X"9D3", X"9D4", X"9D5", 
X"9D5", X"9D6", X"9D7", X"9D8", X"9D9", X"9D9", X"9DA", X"9DB", 
X"9DC", X"9DD", X"9DE", X"9DF", X"9E0", X"9E1", X"9E2", X"9E3", 
X"9E3", X"9E5", X"9E6", X"9E7", X"9E8", X"9E9", X"9EA", X"9EB", 
X"9ED", X"9EE", X"9EF", X"9F0", X"9F2", X"9F3", X"9F4", X"9F6", 
X"9F7", X"9F9", X"9FA", X"9FC", X"9FD", X"9FF", X"A01", X"A02", 
X"A04", X"A06", X"A08", X"A0A", X"A0C", X"A0E", X"A10", X"A12", 
X"A14", X"A16", X"A18", X"A1A", X"A1D", X"A1F", X"A22", X"A24", 
X"A26", X"A29", X"A2C", X"A2E", X"A31", X"A34", X"A37", X"A39", 
X"A3C", X"A3F", X"A43", X"A46", X"A49", X"A4C", X"A4F", X"A53", 
X"A56", X"A5A", X"A5D", X"A61", X"A64", X"A68", X"A6C", X"A70", 
X"A74", X"A78", X"A7C", X"A81", X"A85", X"A89", X"A8D", X"A92", 
X"A97", X"A9B", X"AA0", X"AA4", X"AA9", X"AAE", X"AB3", X"AB8", 
X"ABD", X"AC3", X"AC8", X"ACD", X"AD3", X"AD8", X"ADE", X"AE3", 
X"AE9", X"AEF", X"AF5", X"AFB", X"B01", X"B07", X"B0D", X"B13", 
X"B1A", X"B20", X"B27", X"B2D", X"B34", X"B3B", X"B42", X"B48", 
X"B50", X"B57", X"B5E", X"B65", X"B6C", X"B74", X"B7C", X"B83", 
X"B8B", X"B92", X"B9A", X"BA3", X"BAA", X"BB2", X"BBA", X"BC3", 
X"BCB", X"BD3", X"BDC", X"BE4", X"BEC", X"BF5", X"BFE", X"C07", 
X"C10", X"C19", X"C22", X"C2B", X"C35", X"C3D", X"C47", X"C50", 
X"C5A", X"C63", X"C6D", X"C77", X"C81", X"C8B", X"C94", X"C9E", 
X"CA9", X"CB3", X"CBD", X"CC7", X"CD2", X"CDC", X"CE6", X"CF1", 
X"CFC", X"D06", X"D10", X"D1B", X"D26", X"D32", X"D3D", X"D47", 
X"D52", X"D5E", X"D69", X"D74", X"D7F", X"D8B", X"D96", X"DA1", 
X"DAD", X"DB9", X"DC5", X"DD1", X"DDB", X"DE7", X"DF4", X"E00", 
X"E0B", X"E17", X"E23", X"E2F", X"E3B", X"E47", X"E53", X"E60", 
X"E6B", X"E78", X"E84", X"E91", X"E9D", X"EA9", X"EB6", X"EC2", 
X"ECF", X"EDB", X"EE8", X"EF4", X"F01", X"F0D", X"F1A", X"F27", 
X"F34", X"F41", X"F4C", X"F59", X"F66", X"F73", X"F7F", X"F8C", 
X"F99", X"FA6", X"FB2", X"FBF", X"FCC", X"FD9", X"FE5", X"FF2" 
);

signal data : std_logic_vector(31 downto 0);
signal unsignedIndex : unsigned(11 downto 0) := X"000";

begin

rom_select: process (clk, en)
begin
	if (rising_edge(clk)) then
    if (en = '1') then
		unsignedIndex <= unsigned(address_reg);
		data <= (SIN_ROM(to_integer(unsignedIndex)) & x"00000");
		sin_out <= std_logic_vector(shift_right(signed(data), 20));
    end if;
  end if;
end process rom_select;

end rtl;
