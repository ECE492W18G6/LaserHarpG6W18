----------------------------------------------------------------------------------------------------------
-- Original Authors : Oliver Rarog					                                                    --
-- Date created: March 7, 2018											                                --
--														 	                                            --
-- This component is adapted from the sin_lut component also included in this project, see that         --
-- component for its original and aditional authors.                                 					--
--			                                                                                            --
-- This component takes as an input an index in the range of 0 - 4095 and returns the value at that     --
-- index inside this piano envelope LUT. In order for the output to not be 0, you must enable           --
-- en to '1'.                                                                                       	--
----------------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.all;

entity PianoEnvelope_lut is 

	port(
	-- system signals
	clk 		: in std_logic:= '0'; 
	reset 		: in std_logic:= '0'; 
	en			: in std_logic:= '0';  
	
	-- Current value of the envelope
	index		: in std_logic_vector(11 downto 0);
	data_out 	: out std_logic_vector(31 downto 0)
	);
	
end PianoEnvelope_lut;

architecture rtl of PianoEnvelope_lut is

type rom_type is array (0 to 4095) of std_logic_vector (31 downto 0);

constant ENVELOPE_ROM : rom_type := 
(
X"3f613317", X"3f65d77a", X"3f66afd9", X"3f66458d", X"3f663a02", X"3f64f48a", X"3f654ebe", X"3f684db9", 
X"3f66fa82", X"3f64f0f1", X"3f64ddb7", X"3f65de23", X"3f67cadd", X"3f685f09", X"3f677d8f", X"3f673df3", 
X"3f675601", X"3f6a8538", X"3f6c3873", X"3f6b4899", X"3f69eec6", X"3f695833", X"3f697aeb", X"3f6c75ee", 
X"3f6c137c", X"3f6b65b2", X"3f6a9482", X"3f69f840", X"3f6adf28", X"3f6d4fa2", X"3f6c117a", X"3f6b752d", 
X"3f6accf8", X"3f6d0d32", X"3f709657", X"3f716296", X"3f723924", X"3f73185b", X"3f73ea34", X"3f758ed3", 
X"3f798c0f", X"3f792482", X"3f79ef66", X"3f7b03d2", X"3f7904de", X"3f7c93d9", X"3f7cd0bf", X"3f7d5bc1", 
X"3f7cb93b", X"3f7a17bf", X"3f7b4c2c", X"3f7cd19b", X"3f7c4962", X"3f7c7682", X"3f7a36a3", X"3f781d5c", 
X"3f7b713e", X"3f7a3e8d", X"3f7a7d3e", X"3f79981b", X"3f795420", X"3f791007", X"3f77c0ba", X"3f7663a0", 
X"3f7679c2", X"3f76a1cd", X"3f750d6f", X"3f77f965", X"3f76f3e7", X"3f7655bb", X"3f75c7a9", X"3f773302", 
X"3f791cba", X"3f794d4b", X"3f787beb", X"3f786a9a", X"3f79469d", X"3f7848e9", X"3f7a6d49", X"3f79f5ec", 
X"3f78fa20", X"3f76f561", X"3f76e574", X"3f7a58f4", X"3f79bf84", X"3f79e240", X"3f790661", X"3f7a6bec", 
X"3f790aeb", X"3f7b2977", X"3f7a7839", X"3f7a7dc3", X"3f7addee", X"3f780291", X"3f7b1e06", X"3f7a5c35", 
X"3f7a9266", X"3f788fc6", X"3f7a1b5c", X"3f7b6ada", X"3f7c184e", X"3f7baafb", X"3f7a9ffb", X"3f7b94fd", 
X"3f776b69", X"3f7aa2a1", X"3f79cbb2", X"3f798bb5", X"3f772789", X"3f77f849", X"3f7aa176", X"3f7ad59c", 
X"3f7a5844", X"3f78dd8a", X"3f7ac07c", X"3f785ac6", X"3f7b7af5", X"3f7ada64", X"3f7ac159", X"3f7a15c5", 
X"3f79147e", X"3f7bd5f7", X"3f7acf26", X"3f7b0324", X"3f76df13", X"3f7a42d8", X"3f79585f", X"3f7b7aab", 
X"3f7ae29d", X"3f7a9119", X"3f7ab8aa", X"3f784bc1", X"3f7c782e", X"3f7bf640", X"3f7c48c9", X"3f78b18f", 
X"3f7adc88", X"3f7c9795", X"3f7dc4a4", X"3f7dfa8c", X"3f7bf2dd", X"3f7d91ad", X"3f7aae17", X"3f7ee1a5", 
X"3f7e6b19", X"3f7f1263", X"3f7bdf6b", X"3f7c361e", X"3f7e795e", X"3f7e4002", X"3f7ebd26", X"3f7bb7e9", 
X"3f7e508c", X"3f7bc40f", X"3f7e930a", X"3f7e49bc", X"3f7e5e40", X"3f7d15ea", X"3f7bc885", X"3f7f118a", 
X"3f7e6c26", X"3f7f53bd", X"3f7c238a", X"3f7e63fd", X"3f7e2667", X"3f7f8fa6", X"3f7ff8e8", X"3f7e4144", 
X"3f7e5b9c", X"3f7bbdb6", X"3f7f97f9", X"3f7f43f2", X"3f7ffa17", X"3f7c2b02", X"3f7cd3f0", X"3f7d9a69", 
X"3f7e0af3", X"3f7e7f81", X"3f7bcc0e", X"3f7d2e85", X"3f7a6341", X"3f7dc413", X"3f7d7531", X"3f7da5e5", 
X"3f7a6cbe", X"3f7a0c7b", X"3f7c632f", X"3f7c2f60", X"3f7cd7da", X"3f792b15", X"3f7ab8fb", X"3f78cdf3", 
X"3f7aa84d", X"3f7ad5d3", X"3f798c0c", X"3f77a15b", X"3f748db3", X"3f776242", X"3f76d6af", X"3f774d47", 
X"3f72f8c6", X"3f73883c", X"3f7207fe", X"3f727a6b", X"3f727dd6", X"3f705639", X"3f6fe4db", X"3f6bed1d", 
X"3f6f1d55", X"3f6e41be", X"3f6e5de1", X"3f6aacbb", X"3f6a541c", X"3f6b357b", X"3f6ab5b6", X"3f6b8852", 
X"3f688ae4", X"3f69b981", X"3f67531d", X"3f6a011d", X"3f69b53f", X"3f6913d7", X"3f670d53", X"3f653980", 
X"3f685dd6", X"3f679168", X"3f682bc3", X"3f64ba38", X"3f66509b", X"3f64c56b", X"3f663ba1", X"3f6670f4", 
X"3f653959", X"3f64290a", X"3f610aa4", X"3f64694f", X"3f63b352", X"3f63cdcb", X"3f60767d", X"3f60fa28", 
X"3f614ab9", X"3f61964d", X"3f620818", X"3f5ffe6e", X"3f60f968", X"3f5df94f", X"3f610c2e", X"3f60b19e", 
X"3f609723", X"3f5e0d8c", X"3f5d5851", X"3f5fdbd5", X"3f5f38e5", X"3f5fea92", X"3f5d6d1b", X"3f5eea97", 
X"3f5d630e", X"3f603d6e", X"3f6047bd", X"3f5fcc91", X"3f5ef6c2", X"3f5ddb86", X"3f616429", X"3f60d5ca", 
X"3f619b57", X"3f5f32f0", X"3f60f40d", X"3f60d872", X"3f6274ba", X"3f6344c1", X"3f625bf5", X"3f62a787", 
X"3f607d41", X"3f641c3a", X"3f63fa7b", X"3f648a61", X"3f626b14", X"3f62c743", X"3f64b854", X"3f64bda5", 
X"3f657634", X"3f63936c", X"3f6479ed", X"3f61b800", X"3f650207", X"3f652525", X"3f651081", X"3f6343da", 
X"3f626de4", X"3f64bfbf", X"3f64944a", X"3f652fdc", X"3f62f146", X"3f648342", X"3f633e02", X"3f6509d2", 
X"3f658f26", X"3f64f969", X"3f647fbd", X"3f62ef1b", X"3f660409", X"3f663547", X"3f66cd9e", X"3f64e101", 
X"3f65cf2f", X"3f66357b", X"3f6740b6", X"3f67e7cc", X"3f66b97e", X"3f667366", X"3f642e45", X"3f6719f0", 
X"3f67a8aa", X"3f67db6d", X"3f65b552", X"3f6577d1", X"3f661657", X"3f66ede0", X"3f6781af", X"3f65c7b1", 
X"3f66539b", X"3f63c182", X"3f6609fa", X"3f663f26", X"3f65f38b", X"3f63dde8", X"3f629b6f", X"3f63deb2", 
X"3f643b00", X"3f648f48", X"3f6290d5", X"3f630dbb", X"3f617381", X"3f62b098", X"3f62c856", X"3f6217d7", 
X"3f60d977", X"3f5e92c5", X"3f60de82", X"3f60e249", X"3f6122be", X"3f5eec9f", X"3f5f674b", X"3f5de24e", 
X"3f5ec6ee", X"3f5eda99", X"3f5dc75e", X"3f5d772c", X"3f5afd21", X"3f5cf80a", X"3f5cfa33", X"3f5cf26e", 
X"3f5a5f1b", X"3f59cdec", X"3f5a0082", X"3f5af687", X"3f5b34e5", X"3f598d1b", X"3f59bf34", X"3f57a735", 
X"3f592649", X"3f5912c2", X"3f58b6ae", X"3f567d74", X"3f54d8c3", X"3f561e20", X"3f568d20", X"3f56a7fe", 
X"3f54c86d", X"3f55213e", X"3f53068c", X"3f5412c6", X"3f5401cf", X"3f5389d8", X"3f5218b7", X"3f50b0be", 
X"3f51ecd3", X"3f51ee7b", X"3f520fa2", X"3f4fcc35", X"3f50747a", X"3f4f5b5f", X"3f50c0a7", X"3f50a71b", 
X"3f501a4b", X"3f4fa489", X"3f4e3456", X"3f4f7211", X"3f4f50dc", X"3f4f64d1", X"3f4d355c", X"3f4d1ad9", 
X"3f4d2824", X"3f4e2c39", X"3f4e540a", X"3f4cfb9a", X"3f4d2247", X"3f4bb8ba", X"3f4d4632", X"3f4cf071", 
X"3f4cf83b", X"3f4b08fa", X"3f4ab624", X"3f4b4bdf", X"3f4bf9dc", X"3f4c62e3", X"3f4a3e5d", X"3f4b1932", 
X"3f4a1add", X"3f4c228b", X"3f4c255b", X"3f4bf44a", X"3f4a6b8e", X"3f49f6d6", X"3f4af5b3", X"3f4b2cc0", 
X"3f4b9c3a", X"3f497b79", X"3f49fe33", X"3f48e027", X"3f4aaa5f", X"3f4adb38", X"3f49b66c", X"3f48ed2e", 
X"3f47e854", X"3f4945d1", X"3f490c43", X"3f49736f", X"3f46eeb9", X"3f470a06", X"3f46ab1a", X"3f47c8a6", 
X"3f4811d1", X"3f469d08", X"3f46b2d5", X"3f4566d2", X"3f4780e3", X"3f473ff3", X"3f473d49", X"3f44fdf3", 
X"3f4564b8", X"3f45dd95", X"3f465f86", X"3f46dfa4", X"3f44d473", X"3f45789f", X"3f43bd21", X"3f45dacd", 
X"3f45dd26", X"3f455166", X"3f43c3f8", X"3f439140", X"3f44fc15", X"3f44e475", X"3f457f6e", X"3f42fdb2", 
X"3f43eb70", X"3f42fedb", X"3f44da71", X"3f44ff72", X"3f44168a", X"3f436c59", X"3f4215a5", X"3f440ae9", 
X"3f439ac3", X"3f43dd3b", X"3f40d306", X"3f41d0cf", X"3f413e8f", X"3f42035f", X"3f427b30", X"3f410b9f", 
X"3f40def4", X"3f3ed2af", X"3f40e089", X"3f408640", X"3f4064e9", X"3f3dce1c", X"3f3e5a8a", X"3f3ef6a9", 
X"3f3e915d", X"3f3f2cde", X"3f3d0db5", X"3f3e020e", X"3f3c111f", X"3f3ddde3", X"3f3dd8df", X"3f3d8b4f", 
X"3f3c082b", X"3f3b9919", X"3f3d7068", X"3f3cce01", X"3f3d5023", X"3f3ab143", X"3f3c38cf", X"3f3b0d53", 
X"3f3c4879", X"3f3cec47", X"3f3c1937", X"3f3b8893", X"3f39e7b4", X"3f3c2051", X"3f3bcd0c", X"3f3c058c", 
X"3f38fff1", X"3f3a0883", X"3f39fa16", X"3f3a3711", X"3f3b088b", X"3f39341d", X"3f3995e9", X"3f375166", 
X"3f398cd1", X"3f398abe", X"3f398143", X"3f36cdc2", X"3f36edde", X"3f37e1ae", X"3f376f76", X"3f383671", 
X"3f358db1", X"3f36f741", X"3f34aea7", X"3f367e6b", X"3f3704b9", X"3f36b8c0", X"3f355bac", X"3f34a39d", 
X"3f36708e", X"3f361c16", X"3f36b381", X"3f33d43f", X"3f356d75", X"3f348ad0", X"3f356e06", X"3f36493e", 
X"3f3549ce", X"3f353dbd", X"3f333452", X"3f35fb7e", X"3f35f0ed", X"3f3660eb", X"3f33c15b", X"3f34b14a", 
X"3f350797", X"3f35697d", X"3f365375", X"3f346bd9", X"3f3566b4", X"3f332244", X"3f35b45c", X"3f36130f", 
X"3f362c1d", X"3f341581", X"3f33b94c", X"3f3500b7", X"3f351428", X"3f35f9e2", X"3f335a24", X"3f34e382", 
X"3f32f6e1", X"3f347ff6", X"3f350dce", X"3f34a440", X"3f3397b7", X"3f31c700", X"3f340801", X"3f33efcf", 
X"3f34a945", X"3f321ad5", X"3f338e7d", X"3f328356", X"3f334f29", X"3f342709", X"3f32e9fd", X"3f3338b2", 
X"3f30e9bc", X"3f339392", X"3f339338", X"3f341197", X"3f31ac1a", X"3f322e01", X"3f32508e", X"3f32b380", 
X"3f33a2e8", X"3f319ec8", X"3f32e476", X"3f309568", X"3f32b98d", X"3f32e3da", X"3f32e0ff", X"3f310e95", 
X"3f3000b9", X"3f3199cf", X"3f3185fe", X"3f3267be", X"3f30049f", X"3f319237", X"3f2fb6f6", X"3f312b43", 
X"3f31b1bc", X"3f30f35b", X"3f307a9a", X"3f2e4136", X"3f3054a9", X"3f30129e", X"3f30b412", X"3f2e3f84", 
X"3f2f5c3b", X"3f2e298e", X"3f2f1132", X"3f2fd594", X"3f2e82ad", X"3f2f2977", X"3f2cabdc", X"3f2eef9d", 
X"3f2ed0e2", X"3f2f0f6e", X"3f2d2855", X"3f2d099c", X"3f2d33e1", X"3f2d5ab5", X"3f2e2510", X"3f2c3779", 
X"3f2db5f8", X"3f2b6014", X"3f2d4232", X"3f2d764c", X"3f2d3ec2", X"3f2c6987", X"3f2b4165", X"3f2c58b0", 
X"3f2c37fc", X"3f2ce90d", X"3f2aa060", X"3f2c491b", X"3f2a7878", X"3f2c1528", X"3f2c8192", X"3f2bd3c4", 
X"3f2be44a", X"3f29e138", X"3f2b7153", X"3f2b3ddd", X"3f2b9a58", X"3f299263", X"3f2a615d", X"3f294d6f", 
X"3f2a1f50", X"3f2aa683", X"3f2933ef", X"3f2a0967", X"3f278df2", X"3f2987c5", X"3f2960e5", X"3f2984ce", 
X"3f283b4e", X"3f2806f4", X"3f27d787", X"3f282c42", X"3f28b89c", X"3f26c2e5", X"3f28346e", X"3f25dccb", 
X"3f27cc40", X"3f27d06b", X"3f27a48f", X"3f26e8dc", X"3f25ce89", X"3f268c41", X"3f26a7f8", X"3f271d19", 
X"3f252688", X"3f2654ef", X"3f245f33", X"3f25d2fc", X"3f261c70", X"3f25309b", X"3f2539f0", X"3f23204c", 
X"3f24a424", X"3f2488c7", X"3f24fed5", X"3f234d8a", X"3f23cda3", X"3f22bd41", X"3f23bfdb", X"3f244312", 
X"3f22af87", X"3f235e6d", X"3f2111ea", X"3f231251", X"3f22fe2b", X"3f2321b0", X"3f2187b1", X"3f21356e", 
X"3f20ee7e", X"3f2191e4", X"3f220fc7", X"3f2032a6", X"3f2110ac", X"3f1e85cd", X"3f20570b", X"3f2074d8", 
X"3f1ff95a", X"3f1f0e4a", X"3f1dfc6b", X"3f1e9c18", X"3f1ecbda", X"3f1f4776", X"3f1d6a8d", X"3f1e36a6", 
X"3f1c54e4", X"3f1df6aa", X"3f1e3697", X"3f1d2a8c", X"3f1d2c6b", X"3f1b5905", X"3f1cc340", X"3f1cc4d8", 
X"3f1d1ca7", X"3f1b26c1", X"3f1ba05f", X"3f1a3cbc", X"3f1b9f70", X"3f1bfa2e", X"3f1aab0c", X"3f1b268a", 
X"3f18de46", X"3f1aad69", X"3f1a9f61", X"3f1a888e", X"3f192818", X"3f18edb0", X"3f186b29", X"3f192310", 
X"3f1981ef", X"3f17eb48", X"3f189e99", X"3f16566c", X"3f182e28", X"3f182dba", X"3f17ac40", X"3f16f5af", 
X"3f15df51", X"3f166672", X"3f168111", X"3f16de82", X"3f153129", X"3f1600ef", X"3f13c80b", X"3f1567a6", 
X"3f157978", X"3f14c2c0", X"3f14b938", X"3f12fd2e", X"3f141de4", X"3f13f86f", X"3f14076a", X"3f127e27", 
X"3f12f072", X"3f1178eb", X"3f129c3f", X"3f12c092", X"3f11bb65", X"3f12332c", X"3f1003b0", X"3f11a0a7", 
X"3f116399", X"3f1156eb", X"3f103915", X"3f101030", X"3f0fa5e4", X"3f10276b", X"3f105d09", X"3f0f0564", 
X"3f0fcefc", X"3f0d48f9", X"3f0f37c0", X"3f0f0ae1", X"3f0eb8b7", X"3f0e01df", X"3f0d2ff7", X"3f0d988c", 
X"3f0dbd74", X"3f0ded67", X"3f0c50e6", X"3f0d1b4e", X"3f0aeb0d", X"3f0c6d59", X"3f0c5364", X"3f0bc4e8", 
X"3f0bb206", X"3f09f4aa", X"3f0b246c", X"3f0adfb4", X"3f0b1798", X"3f09bfc6", X"3f0a4a4a", X"3f0916dd", 
X"3f0a2c6c", X"3f0a4d99", X"3f0945c2", X"3f09cf29", X"3f078db2", X"3f09ac78", X"3f096d15", X"3f098eb9", 
X"3f08963c", X"3f089069", X"3f083f03", X"3f08e97a", X"3f093c13", X"3f07d17c", X"3f08a8ab", X"3f067913", 
X"3f08712f", X"3f0848ab", X"3f080efa", X"3f07760d", X"3f06ad14", X"3f075d48", X"3f0774d6", X"3f07e468", 
X"3f067279", X"3f074654", X"3f0589c2", X"3f0743f2", X"3f0745ce", X"3f068bf0", X"3f068a6e", X"3f04dd1d", 
X"3f06847d", X"3f064c13", X"3f06acaf", X"3f054a59", X"3f05bf51", X"3f04809f", X"3f05ba05", X"3f05f31a", 
X"3f04e853", X"3f055a12", X"3f0353dc", X"3f054934", X"3f050696", X"3f051f02", X"3f04151d", X"3f03ee67", 
X"3f03c43e", X"3f0448cf", X"3f04c097", X"3f0392be", X"3f04588f", X"3f0263a2", X"3f0482e5", X"3f0468dc", 
X"3f041b87", X"3f039612", X"3f02bb43", X"3f03c06a", X"3f03ca5b", X"3f045db0", X"3f02f6ad", X"3f03c521", 
X"3f01e8be", X"3f03aca5", X"3f03c928", X"3f032437", X"3f0319ec", X"3f015e54", X"3f02f259", X"3f02916b", 
X"3f02e38c", X"3f016b6d", X"3f01c361", X"3f0088f2", X"3f017ee4", X"3f01d5e0", X"3f00f2c5", X"3f013d88", 
X"3efe3ed7", X"3f010e26", X"3f00c771", X"3f00c77e", X"3eff6f8e", X"3efef47a", X"3efee6c3", X"3eff4d84", 
X"3f002d55", X"3efdc3e7", X"3eff40ae", X"3efa9a8f", X"3efeab98", X"3efe66dd", X"3efdfb9a", X"3efcda33", 
X"3efb0d41", X"3efca655", X"3efc4df3", X"3efd1354", X"3efa62f5", X"3efbb7a0", X"3ef83672", X"3efb4038", 
X"3efb9a3b", X"3efaa0e9", X"3efa77d7", X"3ef70396", X"3efa13e1", X"3ef974a4", X"3ef9efbf", X"3ef778f2", 
X"3ef83b76", X"3ef668c6", X"3ef7d7c4", X"3ef8a568", X"3ef6a6aa", X"3ef75e66", X"3ef2a527", X"3ef67978", 
X"3ef5ee24", X"3ef64179", X"3ef4049f", X"3ef35146", X"3ef2d205", X"3ef2fafb", X"3ef3e867", X"3ef151d7", 
X"3ef283f7", X"3eedc4b8", X"3ef12b4f", X"3ef0d8d1", X"3ef08549", X"3eef3850", X"3eecf389", X"3eee533f", 
X"3eedd640", X"3eeebeab", X"3eec40cc", X"3eed6bdd", X"3eea1c6b", X"3eec444f", X"3eecacb4", X"3eeb7991", 
X"3eeb60c5", X"3ee7853b", X"3eea989c", X"3ee9edee", X"3eeac9aa", X"3ee85532", X"3ee8dc5d", X"3ee7174e", 
X"3ee82c8c", X"3ee9103b", X"3ee71f3e", X"3ee7cff7", X"3ee334ca", X"3ee6a8c4", X"3ee62f9a", X"3ee67fc1", 
X"3ee45cc2", X"3ee37b2c", X"3ee37344", X"3ee3c9e4", X"3ee4f303", X"3ee2cb8d", X"3ee3f57c", X"3edfc04f", 
X"3ee2c556", X"3ee2c2a1", X"3ee24711", X"3ee12a11", X"3ede72ce", X"3ee06433", X"3edff15b", X"3ee11e64", 
X"3ede9668", X"3edf85a0", X"3edc4eda", X"3ede73bb", X"3edef6f0", X"3eddda0c", X"3edd9b80", X"3ed9e450", 
X"3edcbbf9", X"3edbf307", X"3edcd8bf", X"3edaa210", X"3edae452", X"3ed934fe", X"3eda19de", X"3edb2c63", 
X"3ed9a512", X"3eda5ed3", X"3ed68647", X"3ed9a0b0", X"3ed94d56", X"3ed986c4", X"3ed7eac3", X"3ed6ddb5", 
X"3ed754c4", X"3ed7649c", X"3ed8c654", X"3ed6b95a", X"3ed7e32d", X"3ed45921", X"3ed75d59", X"3ed78739", 
X"3ed7240e", X"3ed64675", X"3ed3c4ca", X"3ed5f00b", X"3ed569eb", X"3ed68d66", X"3ed42f07", X"3ed4f051", 
X"3ed21624", X"3ed3fd56", X"3ed4b7d3", X"3ed3cd7c", X"3ed3a171", X"3ed04bdc", X"3ed3035d", X"3ed25b65", 
X"3ed3048e", X"3ed101d9", X"3ed0cac0", X"3ecfb0fe", X"3ed05565", X"3ed17972", X"3ecfdd76", X"3ed07c37", 
X"3ecc9d2a", X"3ecfaaa9", X"3ecf5ea0", X"3ecfb4f2", X"3ece60b7", X"3ecce982", X"3ecd7573", X"3ecd6956", 
X"3ece9d36", X"3eccc05b", X"3ecd9c4d", X"3eca2384", X"3eccea96", X"3ecd2f1b", X"3eccd633", X"3ecc4726", 
X"3ec9eb62", X"3ecbb9f3", X"3ecb3300", X"3ecc4d34", X"3eca6204", X"3ecad652", X"3ec8c14c", X"3eca3b4c", 
X"3ecb1caa", X"3eca15d1", X"3eca07c3", X"3ec6b637", X"3ec96b88", X"3ec8ff32", X"3ec9c7c9", X"3ec81eff", 
X"3ec7a058", X"3ec6a789", X"3ec723b3", X"3ec82dba", X"3ec68e24", X"3ec6f9ea", X"3ec32525", X"3ec5e2ef", 
X"3ec5a250", X"3ec5f02c", X"3ec4ae07", X"3ec33179", X"3ec351da", X"3ec336c4", X"3ec471db", X"3ec2e1c0", 
X"3ec36a81", X"3ec05aa5", X"3ec28532", X"3ec2dc77", X"3ec27765", X"3ec1e2c9", X"3ebf625d", X"3ec12e2e", 
X"3ec0dba8", X"3ec214ec", X"3ec0881b", X"3ec0afa0", X"3ebe9aa3", X"3ec01a8a", X"3ec0ea95", X"3ebfeb95", 
X"3ebfd5b7", X"3ebc9880", X"3ebef304", X"3ebe9fba", X"3ebf724b", X"3ebe0194", X"3ebd59c1", X"3ebc2359", 
X"3ebcd750", X"3ebdeed0", X"3ebcb525", X"3ebd036c", X"3eb98237", X"3ebbe7db", X"3ebbcf3b", X"3ebbe113", 
X"3ebacbf8", X"3eb92db1", X"3eb9a9fc", X"3eb9b91e", X"3ebaf02a", X"3eb986d6", X"3eb9cc37", X"3eb6f28e", 
X"3eb8f2a5", X"3eb93e98", X"3eb8d425", X"3eb84c30", X"3eb5d701", X"3eb760fe", X"3eb70921", X"3eb811f0", 
X"3eb69e11", X"3eb6a528", X"3eb48768", X"3eb5f9ba", X"3eb6ae7e", X"3eb603cb", X"3eb5fc5c", X"3eb32159", 
X"3eb562cb", X"3eb52334", X"3eb5a6c2", X"3eb468ae", X"3eb3b566", X"3eb322ae", X"3eb3e77e", X"3eb4f8e3", 
X"3eb3ea37", X"3eb421ac", X"3eb116fa", X"3eb35f4d", X"3eb3455a", X"3eb368b3", X"3eb2906e", X"3eb0fac2", 
X"3eb14617", X"3eb14545", X"3eb25789", X"3eb11ec8", X"3eb15ead", X"3eae82b3", X"3eb06042", X"3eb077f8", 
X"3eb052b3", X"3eafe017", X"3eadcd88", X"3eaf36b7", X"3eaee940", X"3eafbbd2", X"3eae94a9", X"3eae7c9c", 
X"3eacaa3e", X"3eadf5af", X"3eae9bae", X"3eae0b23", X"3eadea8f", X"3eab42f6", X"3ead3864", X"3eacc8c4", 
X"3ead6ea6", X"3eac66e9", X"3eaba6a9", X"3eaad0a4", X"3eab7cfc", X"3eac7043", X"3eab7658", X"3eaba1c3", 
X"3ea8c338", X"3eab13b0", X"3eaae27c", X"3eab2933", X"3eaa44b1", X"3ea90fe9", X"3ea98109", X"3ea9ac3c", 
X"3eaab984", X"3ea9ac95", X"3ea9d87d", X"3ea75829", X"3ea95213", X"3ea99a27", X"3ea96db5", X"3ea8cde2", 
X"3ea6bdd6", X"3ea80864", X"3ea7d762", X"3ea8d265", X"3ea7b75a", X"3ea77a14", X"3ea58cf6", X"3ea6fa25", 
X"3ea785ee", X"3ea6d404", X"3ea6a388", X"3ea40bc0", X"3ea607a5", X"3ea5a57f", X"3ea65084", X"3ea5438f", 
X"3ea4afac", X"3ea3e82b", X"3ea4c866", X"3ea5a114", X"3ea4ca4d", X"3ea4d7c3", X"3ea24941", X"3ea49df2", 
X"3ea48b71", X"3ea4aa56", X"3ea3c1ec", X"3ea27a77", X"3ea2e9fb", X"3ea33356", X"3ea459bb", X"3ea3595a", 
X"3ea362e8", X"3ea0f8bf", X"3ea34fae", X"3ea39094", X"3ea35c13", X"3ea2c696", X"3ea0ef67", X"3ea26fd6", 
X"3ea2481e", X"3ea345b0", X"3ea22a82", X"3ea2082e", X"3ea00b64", X"3ea1b9b6", X"3ea26aaf", X"3ea1e277", 
X"3ea1906d", X"3e9f163f", X"3ea11eab", X"3ea0bef7", X"3ea15e83", X"3ea02940", X"3e9f8285", X"3e9e71ac", 
X"3e9f395b", X"3ea03c09", X"3e9f82cc", X"3e9f5131", X"3e9c84b5", X"3e9ec1c9", X"3e9e8447", X"3e9eb74e", 
X"3e9dd639", X"3e9c9bf1", X"3e9cea49", X"3e9ce98e", X"3e9de724", X"3e9cf375", X"3e9d0c7f", X"3e9a7007", 
X"3e9cb2f4", X"3e9cf3fb", X"3e9cd653", X"3e9c35ee", X"3e9a7ddb", X"3e9be4b3", X"3e9ba5a1", X"3e9c8f69", 
X"3e9b70ae", X"3e9b4a2a", X"3e99563d", X"3e9aef71", X"3e9bbc5a", X"3e9b4bbc", X"3e9adf55", X"3e9855f4", 
X"3e9a4c59", X"3e99e827", X"3e9a7b9b", X"3e99671f", X"3e98ce96", X"3e97bc36", X"3e9847a0", X"3e993b9f", 
X"3e987b97", X"3e98551b", X"3e954675", X"3e977d94", X"3e975043", X"3e979b8b", X"3e9690ca", X"3e958335", 
X"3e959328", X"3e957d1e", X"3e9675d1", X"3e958fdb", X"3e95a384", X"3e92fa32", X"3e94e233", X"3e952701", 
X"3e951639", X"3e945d94", X"3e92a213", X"3e93e409", X"3e9398c5", X"3e946a71", X"3e937edc", X"3e9388c1", 
X"3e91c7dc", X"3e932244", X"3e93dad7", X"3e936d9b", X"3e9330b5", X"3e90ade4", X"3e92d37a", X"3e929c59", 
X"3e933306", X"3e922aac", X"3e91db5c", X"3e910b43", X"3e91c11e", X"3e92abae", X"3e920381", X"3e91fb69", 
X"3e8f27f9", X"3e9171cc", X"3e91860c", X"3e91bb1e", X"3e90c639", X"3e8f923b", X"3e8fc295", X"3e8fd222", 
X"3e90c0a6", X"3e8ff5e2", X"3e90051b", X"3e8d7a77", X"3e8f3e93", X"3e8f8e25", X"3e8f7cdd", X"3e8eda6f", 
X"3e8cf57f", X"3e8e3b0d", X"3e8e15ca", X"3e8ee10f", X"3e8df16f", X"3e8dfd3b", X"3e8c45d0", X"3e8d955f", 
X"3e8e30d8", X"3e8dea0c", X"3e8d9c40", X"3e8b2766", X"3e8d2352", X"3e8d0909", X"3e8d8eaf", X"3e8c87ce", 
X"3e8c03b7", X"3e8b4064", X"3e8c0221", X"3e8cdab2", X"3e8c5ad9", X"3e8c4dd7", X"3e89bcc0", X"3e8bc3b8", 
X"3e8bc6fc", X"3e8c091a", X"3e8b25ac", X"3e89d57e", X"3e8a267a", X"3e8a6cea", X"3e8b55dd", X"3e8a7866", 
X"3e8a8b4a", X"3e8808c4", X"3e89d932", X"3e8a2b26", X"3e8a395e", X"3e899791", X"3e879853", X"3e88db6c", 
X"3e88cfbc", X"3e898fd9", X"3e88886c", X"3e886572", X"3e8674bc", X"3e87dac2", X"3e8873e6", X"3e883d83", 
X"3e87ec97", X"3e857415", X"3e871f70", X"3e870083", X"3e8780f0", X"3e869b01", X"3e85e3d2", X"3e852d6e", 
X"3e85fea5", X"3e86b6e2", X"3e862ced", X"3e86389d", X"3e83a265", X"3e859208", X"3e859181", X"3e85e309", 
X"3e85295b", X"3e83ec76", X"3e8430f8", X"3e848da2", X"3e85394a", X"3e847f6c", X"3e848b46", X"3e822645", 
X"3e84150e", X"3e844859", X"3e8456e3", X"3e83da4b", X"3e820013", X"3e830275", X"3e82fea5", X"3e839208", 
X"3e82c80a", X"3e828f19", X"3e80d311", X"3e823c85", X"3e829081", X"3e8259b7", X"3e821c65", X"3e7f8d79", 
X"3e816361", X"3e813b0d", X"3e81b111", X"3e80eaf0", X"3e804957", X"3e7e8ef5", X"3e801d57", X"3e808cdc", 
X"3e801ffe", X"3e802039", X"3e7b20bc", X"3e7eae4b", X"3e7e48d2", X"3e7ef0f6", X"3e7d9927", X"3e7b5e15", 
X"3e7aea12", X"3e7ba7de", X"3e7c9e79", X"3e7b88bb", X"3e7b9a1e", X"3e76d32c", X"3e7a4988", X"3e7a376d", 
X"3e7a46ba", X"3e796b2c", X"3e75efb2", X"3e778b9f", X"3e778b20", X"3e788653", X"3e773602", X"3e76f6ab", 
X"3e72d639", X"3e75cd68", X"3e7621c2", X"3e75d804", X"3e7590e6", X"3e70ffea", X"3e73947d", X"3e733941", 
X"3e74218a", X"3e7297b4", X"3e715d21", X"3e6e9958", X"3e7069da", X"3e710d26", X"3e706453", X"3e706626", 
X"3e6b05a4", X"3e6e2a46", X"3e6db121", X"3e6e2b2c", X"3e6cf7a8", X"3e6a964e", X"3e6a0696", X"3e6ae2b5", 
X"3e6ba624", X"3e6aa82b", X"3e6ab8b9", X"3e657310", X"3e68ca81", X"3e68aa5b", X"3e68dc19", X"3e683503", 
X"3e64cd79", X"3e65f5bf", X"3e65f933", X"3e66e32f", X"3e6588ac", X"3e654edd", X"3e611111", X"3e641818", 
X"3e643625", X"3e640fa0", X"3e63bd4a", X"3e5f7b7c", X"3e61e223", X"3e6187d0", X"3e622907", X"3e60b1d5", 
X"3e5fa1ef", X"3e5d32de", X"3e5f4717", X"3e5fcb53", X"3e5f271b", X"3e5f1ac8", X"3e59d758", X"3e5d77d7", 
X"3e5d1bb1", X"3e5d94ca", X"3e5c638f", X"3e5a506c", X"3e5997cf", X"3e5a8529", X"3e5b375e", X"3e5a0e72", 
X"3e5a2bf6", X"3e550b83", X"3e5850d2", X"3e57f0ec", X"3e584188", X"3e5771cc", X"3e549316", X"3e55881a", 
X"3e557b90", X"3e562636", X"3e54e658", X"3e54df87", X"3e5117cc", X"3e53f437", X"3e53e3d5", X"3e53a2d8", 
X"3e534da6", X"3e4f32d0", X"3e51e02f", X"3e517e60", X"3e521d51", X"3e50c7ad", X"3e4fe3b7", X"3e4d7266", 
X"3e4fa63e", X"3e4fdebd", X"3e4f23be", X"3e4f0abc", X"3e4a5642", X"3e4dc53c", X"3e4d227c", X"3e4dac33", 
X"3e4c6938", X"3e4ab50c", X"3e49d7b9", X"3e4a8b3c", X"3e4afad4", X"3e4a0e3a", X"3e4a5084", X"3e458c9d", 
X"3e48a4d5", X"3e483862", X"3e487d17", X"3e47b544", X"3e44d02f", X"3e45c67d", X"3e45ca7f", X"3e4678c0", 
X"3e454b6b", X"3e454158", X"3e414069", X"3e44038a", X"3e43cd3d", X"3e43a6e7", X"3e435601", X"3e3efc67", 
X"3e4169b7", X"3e40fdfe", X"3e41b1d4", X"3e407885", X"3e3fafec", X"3e3d2dca", X"3e3ef885", X"3e3f024e", 
X"3e3e772b", X"3e3e80d4", X"3e3a207f", X"3e3d417a", X"3e3c97c1", X"3e3d0f2b", X"3e3c0165", X"3e3a5b6c", 
X"3e39cd21", X"3e3a7f1f", X"3e3b0609", X"3e3a29c4", X"3e3a75d9", X"3e3604a1", X"3e391801", X"3e38a30a", 
X"3e391244", X"3e387cd2", X"3e357664", X"3e366180", X"3e366142", X"3e372a6d", X"3e3624f2", X"3e360725", 
X"3e321318", X"3e34a556", X"3e347806", X"3e3494a9", X"3e344e19", X"3e305259", X"3e329e5c", X"3e324375", 
X"3e32eb18", X"3e31d119", X"3e311730", X"3e2f1d2f", X"3e30cf94", X"3e30f189", X"3e308ac0", X"3e3092ef", 
X"3e2c8a6a", X"3e2f4262", X"3e2e9fb2", X"3e2f6164", X"3e2e6ddf", X"3e2cbcc5", X"3e2c1d84", X"3e2cc2f0", 
X"3e2d57c5", X"3e2c9e25", X"3e2cd671", X"3e2895db", X"3e2b6537", X"3e2ae9ef", X"3e2b87e4", X"3e2aff59", 
X"3e282cd9", X"3e2902c7", X"3e2923e6", X"3e29d5b1", X"3e2904f9", X"3e28c90a", X"3e25943a", X"3e282609", 
X"3e2803a2", X"3e282f26", X"3e27f5c6", X"3e245da3", X"3e2673de", X"3e260ed8", X"3e26f68e", X"3e25f0c4", 
X"3e25145a", X"3e2335ed", X"3e24add7", X"3e24b769", X"3e24709d", X"3e2478c8", X"3e207cf7", X"3e230aed", 
X"3e224480", X"3e2322e5", X"3e22610e", X"3e20b4e9", X"3e2026f9", X"3e20baed", X"3e211fcb", X"3e20af86", 
X"3e20cc64", X"3e1d2525", X"3e1fc5b2", X"3e1f27b4", X"3e1fbe93", X"3e1f4cb5", X"3e1c9252", X"3e1d6369", 
X"3e1d71e0", X"3e1e1d7c", X"3e1d6ef7", X"3e1d16b1", X"3e1a471d", X"3e1c889f", X"3e1c1252", X"3e1c5702", 
X"3e1c1f2c", X"3e18e5e8", X"3e1af079", X"3e1a4ff9", X"3e1b3358", X"3e1a7765", X"3e19b7b2", X"3e1800cc", 
X"3e193ea4", X"3e192d7d", X"3e1932b8", X"3e193a2f", X"3e15c30b", X"3e1819c0", X"3e175336", X"3e1846c6", 
X"3e17aaae", X"3e15f662", X"3e158f4d", X"3e164c13", X"3e16b196", X"3e167a34", X"3e166e98", X"3e130449", 
X"3e157570", X"3e14acdc", X"3e155c6e", X"3e150a5d", X"3e128b33", X"3e136ac8", X"3e134665", X"3e13fe89", 
X"3e13945e", X"3e135b74", X"3e10b83f", X"3e12a34d", X"3e121c0f", X"3e12a0e0", X"3e1296a8", X"3e0fc779", 
X"3e117400", X"3e10dab7", X"3e11c71f", X"3e1149f1", X"3e1082f5", X"3e0f1206", X"3e107671", X"3e104ec7", 
X"3e1090eb", X"3e109662", X"3e0d73ff", X"3e0f8a4b", X"3e0ec2bf", X"3e0fbf41", X"3e0f6221", X"3e0dc24a", 
X"3e0d5e1e", X"3e0e189e", X"3e0e65d8", X"3e0e5bc5", X"3e0e456c", X"3e0b0708", X"3e0d4f43", X"3e0c756e", 
X"3e0d508d", X"3e0d30df", X"3e0af9fd", X"3e0b882f", X"3e0b7904", X"3e0c1dd5", X"3e0be19c", X"3e0bab37", 
X"3e0979de", X"3e0b36f2", X"3e0a7541", X"3e0b3289", X"3e0b2ce5", X"3e08939c", X"3e09e54f", X"3e093d08", 
X"3e0a23f1", X"3e09ea50", X"3e090a4b", X"3e077c1f", X"3e08d836", X"3e088b4d", X"3e08daf0", X"3e08dacd", 
X"3e05c2ee", X"3e07c4c6", X"3e06f3e4", X"3e07e5c2", X"3e07b181", X"3e0630db", X"3e05cbed", X"3e069024", 
X"3e06a170", X"3e068ce6", X"3e0667ba", X"3e03ccd3", X"3e05dd8c", X"3e04d83a", X"3e05b494", X"3e0574e3", 
X"3e036ef5", X"3e03c21c", X"3e039eda", X"3e041f5c", X"3e041945", X"3e03b9f1", X"3e01683b", X"3e02eb87", 
X"3e021e04", X"3e02d757", X"3e02d284", X"3e0066e1", X"3e01791b", X"3e00cd66", X"3e01a304", X"3e018bec", 
X"3e00ba54", X"3dfe7afe", X"3e008bb9", X"3e0021c7", X"3e008250", X"3e007df0", X"3dfb7e64", X"3dfe94ef", 
X"3dfce8f6", X"3dfe8ecc", X"3dfe1cee", X"3dfb5a8f", X"3dfa3e4f", X"3dfb89d6", X"3dfb3266", X"3dfb96aa", 
X"3dfb3df9", X"3df67739", X"3df9ac05", X"3df792f0", X"3df91c1e", X"3df8f951", X"3df57d46", X"3df5cff3", 
X"3df593db", X"3df67de5", X"3df6b4c9", X"3df60b99", X"3df1764b", X"3df431bb", X"3df2981d", X"3df45a47", 
X"3df473c5", X"3defda6f", X"3df0e613", X"3deff848", X"3df180a4", X"3df18e6c", X"3defe067", X"3dec4178", 
X"3dee9139", X"3ded9779", X"3deeed60", X"3deedeed", X"3de9df6f", X"3debfda8", X"3dea7a23", X"3dec31d1", 
X"3dec41a5", X"3dea0949", X"3de85dd1", X"3de93507", X"3de92990", X"3dea1e13", X"3dea124d", X"3de5bf39", 
X"3de81073", X"3de5d231", X"3de7e21a", X"3de8070f", X"3de50bfd", X"3de4ad17", X"3de47e4a", X"3de54016", 
X"3de5cbfc", X"3de51e89", X"3de10c21", X"3de3b39c", X"3de222f9", X"3de3d74a", X"3de3e0b1", X"3ddff21b", 
X"3de1075b", X"3de08e03", X"3de1d7d9", X"3de237ef", X"3de0b00e", X"3ddda041", X"3ddf9fe0", X"3ddeadbf", 
X"3de01325", X"3de008aa", X"3ddbfa41", X"3dddada8", X"3ddc2153", X"3dddf9c3", X"3dde3c40", X"3ddc4b5b", 
X"3ddaa2ac", X"3ddb74f6", X"3ddaf495", X"3ddc1c59", X"3ddc03b2", X"3dd8529b", X"3dda5be5", X"3dd83cd0", 
X"3dda2c6b", X"3dda5fbc", X"3dd7ecd1", X"3dd716a0", X"3dd71b06", X"3dd764ee", X"3dd84026", X"3dd7a3a2", 
X"3dd46413", X"3dd69ab4", X"3dd4e512", X"3dd686ee", X"3dd69725", X"3dd3763e", X"3dd419fe", X"3dd38368", 
X"3dd48e3a", X"3dd4f869", X"3dd3e700", X"3dd1bcec", X"3dd35d49", X"3dd1b2f6", X"3dd341e6", X"3dd340ee", 
X"3dd01de2", X"3dd1864d", X"3dcfd34f", X"3dd173eb", X"3dd1ccb4", X"3dd05b75", X"3dcec547", X"3dcfad83", 
X"3dcec4f2", X"3dd01aff", X"3dcfe380", X"3dccac64", X"3dce48af", X"3dcc9172", X"3dce9301", X"3dcee7c6", 
X"3dcc53ea", X"3dcb83ca", X"3dcc107b", X"3dcc5078", X"3dcd67d6", X"3dccd9ef", X"3dc9ff1b", X"3dcbd167", 
X"3dc9fbf1", X"3dcc1e3c", X"3dcc622f", X"3dc99ca5", X"3dc99bb1", X"3dc90450", X"3dc9d674", X"3dcaa19a", 
X"3dc9bb1c", X"3dc777e8", X"3dc91d92", X"3dc76afb", X"3dc9526a", X"3dc9795f", X"3dc6e299", X"3dc79062", 
X"3dc63d90", X"3dc7fe8c", X"3dc8962d", X"3dc7288e", X"3dc5a678", X"3dc6c015", X"3dc612e8", X"3dc7d9a3", 
X"3dc7afd4", X"3dc4bc06", X"3dc5d597", X"3dc44c32", X"3dc67836", X"3dc7000a", X"3dc4c829", X"3dc3b987", 
X"3dc44214", X"3dc4260d", X"3dc57648", X"3dc4f0fc", X"3dc25538", X"3dc3ef05", X"3dc1ef17", X"3dc3f7d0", 
X"3dc440b7", X"3dc228a7", X"3dc1e3eb", X"3dc165e5", X"3dc21e89", X"3dc31f11", X"3dc23fc5", X"3dc03656", 
X"3dc1c638", X"3dc027c7", X"3dc2726f", X"3dc29686", X"3dc01e29", X"3dc06448", X"3dbf30f1", X"3dc0a199", 
X"3dc18a5d", X"3dc0115f", X"3dbe1a4c", X"3dbf3cbf", X"3dbe38d4", X"3dc01407", X"3dbff34e", X"3dbd6a8f", 
X"3dbe6244", X"3dbca472", X"3dbe756b", X"3dbf042e", X"3dbd8508", X"3dbc2e77", X"3dbccd26", X"3dbc6997", 
X"3dbe0939", X"3dbda11d", X"3dbb6f4d", X"3dbca706", X"3dba771b", X"3dbcade1", X"3dbd0a6b", X"3dbb4a88", 
X"3dbab9b7", X"3dba5276", X"3dbaa38f", X"3dbc04fd", X"3dbb5431", X"3db96240", X"3dbac9bb", X"3db8cbc6", 
X"3dbae71d", X"3dbb13e3", X"3db9221f", X"3db92ad9", X"3db81dcf", X"3db971e9", X"3dba7219", X"3db94bf4", 
X"3db7543c", X"3db8d263", X"3db78fb9", X"3db9a6de", X"3db9841a", X"3db77991", X"3db81628", X"3db68a3b", 
X"3db8927b", X"3db9344c", X"3db7c310", X"3db650b3", X"3db71a13", X"3db6767c", X"3db86e06", X"3db80d67", 
X"3db5eb49", X"3db719ed", X"3db4f995", X"3db72ff0", X"3db7b468", X"3db63fc2", X"3db5416c", X"3db5201f", 
X"3db5b0e0", X"3db741dc", X"3db6a06a", X"3db4b8bd", X"3db616c8", X"3db4040b", X"3db68700", X"3db6c936", 
X"3db525b2", X"3db4cb4b", X"3db40bc7", X"3db56bb5", X"3db67a85", X"3db58f41", X"3db3e564", X"3db545b5", 
X"3db3bb1c", X"3db5f917", X"3db5ecf4", X"3db46309", X"3db50c91", X"3db37934", X"3db53488", X"3db5f584", 
X"3db4eb82", X"3db398c6", X"3db48025", X"3db40a22", X"3db5c25a", X"3db56f94", X"3db3dd8b", X"3db51572", 
X"3db303c6", X"3db56373", X"3db5d1b1", X"3db4ad3f", X"3db3dde5", X"3db40143", X"3db483f0", X"3db5e553", 
X"3db56065", X"3db38b7d", X"3db509d1", X"3db3284f", X"3db59ea2", X"3db5ce73", X"3db4c358", X"3db48c3a", 
X"3db3a6bb", X"3db50a19", X"3db62e0e", X"3db59001", X"3db3fd67", X"3db53220", X"3db3eb4e", X"3db5ed05", 
X"3db5eb7a", X"3db4c3f6", X"3db5321f", X"3db34695", X"3db54608", X"3db6078a", X"3db55ad3", X"3db43b01", 
X"3db4da77", X"3db43d5b", X"3db5d103", X"3db58f4e", X"3db4521e", X"3db5aff7", X"3db384cd", X"3db593f7", 
X"3db600e8", X"3db54812", X"3db4c2ff", X"3db4a61a", X"3db52f4f", X"3db65ca6", X"3db5c761", X"3db46719", 
X"3db5f04b", X"3db42d8b", X"3db62371", X"3db639bb", X"3db514a1", X"3db50e02", X"3db3dc00", X"3db5670a", 
X"3db66216", X"3db59d82", X"3db3ddf3", X"3db5211b", X"3db3b5e4", X"3db5e9e0", X"3db5bc5c", X"3db45725", 
X"3db4ce85", X"3db2e5d6", X"3db4e3be", X"3db5b563", X"3db4d3b0", X"3db3586d", X"3db3b399", X"3db36934", 
X"3db50e1e", X"3db49f00", X"3db33ad6", X"3db46013", X"3db1fb73", X"3db41fa4", X"3db47bdf", X"3db37abc", 
X"3db2e4ab", X"3db2440c", X"3db2c504", X"3db3fee3", X"3db3622a", X"3db1ddcb", X"3db36e3f", X"3db1654d", 
X"3db37339", X"3db36337", X"3db25d8e", X"3db2a4de", X"3db128d3", X"3db2861a", X"3db36757", X"3db2a9b6", 
X"3db14103", X"3db2475c", X"3db15a74", X"3db31321", X"3db2b1e7", X"3db15bdc", X"3db22211", X"3daffcfb", 
X"3db1f8fc", X"3db277f9", X"3db17abc", X"3db05d1f", X"3db05dad", X"3db093cb", X"3db22882", X"3db193c2", 
X"3dafe2df", X"3db13cec", X"3daf1b07", X"3db15688", X"3db1954b", X"3db0bda3", X"3db02811", X"3daf395c", 
X"3daffa6d", X"3db1395f", X"3db0ae09", X"3daf4512", X"3db0577b", X"3dae9c27", X"3db0534d", X"3db055ec", 
X"3daf8bf6", X"3dafe68c", X"3dae0b6c", X"3daf4160", X"3db00cee", X"3daf7f68", X"3dae7a08", X"3daf4873", 
X"3dae351f", X"3dafaf24", X"3daf54d2", X"3dae3c29", X"3daf52ef", X"3dad3dbc", X"3daebcd7", X"3daf2ebd", 
X"3dae8839", X"3dad7e27", X"3dad5a62", X"3dad5941", X"3daea6d5", X"3dae1208", X"3dac8996", X"3dad9400", 
X"3dab633c", X"3dad54d9", X"3dad88bd", X"3dac90cb", X"3dac0a5e", X"3daacd7c", X"3dab9215", X"3dacb6f9", 
X"3dac0498", X"3daa7093", X"3dab64c9", X"3da9b720", X"3dab88f4", X"3dab545f", X"3daa5996", X"3daaaec5", 
X"3da8bf68", X"3da9ee8a", X"3daaa7df", X"3da9ec4b", X"3da8a6fc", X"3da90033", X"3da8078e", X"3da95522", 
X"3da8d2d0", X"3da7bc9d", X"3da8c61e", X"3da64b74", X"3da7b3d7", X"3da7fb04", X"3da72bf1", X"3da6a144", 
X"3da5f9a4", X"3da5f563", X"3da70ba9", X"3da66d19", X"3da52c79", X"3da6747e", X"3da47f3d", X"3da60739", 
X"3da5e740", X"3da4fc37", X"3da4e8d2", X"3da3776e", X"3da46971", X"3da54594", X"3da47413", X"3da2f619", 
X"3da3b820", X"3da2be5b", X"3da44368", X"3da3cf08", X"3da2b5c4", X"3da346e3", X"3da141c5", X"3da2e058", 
X"3da3703d", X"3da2aa46", X"3da1ade1", X"3da1af83", X"3da154bc", X"3da2bd76", X"3da24764", X"3da1422e", 
X"3da237a3", X"3da04251", X"3da199c4", X"3da1db3e", X"3da1528a", X"3da0f31d", X"3da01a8e", X"3da07439", 
X"3da1816c", X"3da0ecb7", X"3da005e6", X"3da11709", X"3d9f7757", X"3da0cd1b", X"3da0a800", X"3d9ff578", 
X"3da05e64", X"3d9ede74", X"3d9fd8b4", X"3da08c93", X"3d9fdf83", X"3d9ec383", X"3d9f775e", X"3d9e8253", 
X"3d9ffb47", X"3d9f8791", X"3d9e7c86", X"3d9f23cd", X"3d9d66ec", X"3d9ec6a3", X"3d9f51a9", X"3d9e87aa", 
X"3d9dad4a", X"3d9d616d", X"3d9d7678", X"3d9ec833", X"3d9e2987", X"3d9d0174", X"3d9dea50", X"3d9bf824", 
X"3d9dabd0", X"3d9dc1d3", X"3d9d0cc6", X"3d9cf586", X"3d9bd3f7", X"3d9c5ee0", X"3d9d59dd", X"3d9ca66d", 
X"3d9b9ff6", X"3d9c70ac", X"3d9aeb75", X"3d9c524d", X"3d9bfeac", X"3d9b5abc", X"3d9bf1cf", X"3d9a2537", 
X"3d9b0fc0", X"3d9ba428", X"3d9aefd6", X"3d9a5bf1", X"3d9a8876", X"3d99e757", X"3d9b11e0", X"3d9a84a2", 
X"3d99ce1b", X"3d9ae53c", X"3d98ecba", X"3d9a5fc9", X"3d9a8c8f", X"3d99c943", X"3d99898d", X"3d98db27", 
X"3d990a0d", X"3d9a1b22", X"3d9956f7", X"3d98444f", X"3d99500c", X"3d97db6d", X"3d995e2e", X"3d992b5d", 
X"3d9868cc", X"3d988814", X"3d97351e", X"3d983973", X"3d99154c", X"3d984753", X"3d977fee", X"3d98230c", 
X"3d974caf", X"3d98aff3", X"3d9860b0", X"3d97b204", X"3d986de6", X"3d96c180", X"3d97f5e8", X"3d98762b", 
X"3d97e524", X"3d978edd", X"3d979b39", X"3d971d38", X"3d983bfe", X"3d97b2d6", X"3d972af3", X"3d985d5b", 
X"3d96ba4e", X"3d97e31b", X"3d980130", X"3d9765ca", X"3d97850e", X"3d96c2a6", X"3d974262", X"3d982131", 
X"3d9761cb", X"3d96be5b", X"3d97cf69", X"3d967329", X"3d97fd8f", X"3d97c87b", X"3d96e808", X"3d9758e7", 
X"3d961de6", X"3d971d6e", X"3d97e5d7", X"3d96febf", X"3d96309a", X"3d96afb5", X"3d95eca6", X"3d975634", 
X"3d96d4af", X"3d95fa0f", X"3d96c74b", X"3d95033e", X"3d965a01", X"3d96c625", X"3d95f47f", X"3d95bd32", 
X"3d9569e7", X"3d95709b", X"3d9689da", X"3d95d0ac", X"3d951846", X"3d962b5f", X"3d945676", X"3d95afb8", 
X"3d95a83e", X"3d94da57", X"3d953be5", X"3d942297", X"3d9496c5", X"3d956051", X"3d94855f", X"3d93d480", 
X"3d94a754", X"3d937378", X"3d94a200", X"3d944520", X"3d938d8a", X"3d9466d2", X"3d92bf29", X"3d93d352", 
X"3d944b98", X"3d934f50", X"3d92e440", X"3d92fe2b", X"3d92a9fe", X"3d93d19d", X"3d932b5e", X"3d9236c6", 
X"3d93493f", X"3d918e3f", X"3d92ff27", X"3d932a01", X"3d922867", X"3d921043", X"3d916136", X"3d91c79d", 
X"3d92d83c", X"3d920c78", X"3d912684", X"3d92158d", X"3d90b21b", X"3d91f3e8", X"3d91f859", X"3d913af6", 
X"3d9192bf", X"3d90481b", X"3d911235", X"3d91bf35", X"3d90f6d0", X"3d908e9f", X"3d914531", X"3d90494d", 
X"3d915de5", X"3d910597", X"3d905a02", X"3d91726b", X"3d8fdd52", X"3d90cc79", X"3d912ab1", X"3d905797", 
X"3d902298", X"3d90268b", X"3d8feef4", X"3d90d905", X"3d903a5e", X"3d8f720f", X"3d909683", X"3d8f042d", 
X"3d90546a", X"3d908a5e", X"3d8f9572", X"3d8fa40c", X"3d8eec70", X"3d8f7602", X"3d90601e", X"3d8f8db5", 
X"3d8ea9da", X"3d8f9295", X"3d8e2c2e", X"3d8f9d36", X"3d8f7751", X"3d8e7b61", X"3d8efa16", X"3d8d9fb3", 
X"3d8e7343", X"3d8f1d06", X"3d8e31ea", X"3d8dae16", X"3d8e16fd", X"3d8d68e1", X"3d8e72a8", X"3d8dedc6", 
X"3d8d1468", X"3d8e22fc", X"3d8c5c0f", X"3d8d7181", X"3d8dbbb2", X"3d8cd08f", X"3d8cdf82", X"3d8c7c31", 
X"3d8c612f", X"3d8d3054", X"3d8c7702", X"3d8bb05a", X"3d8cda09", X"3d8b3ca1", X"3d8c6019", X"3d8c53e0", 
X"3d8b776b", X"3d8c03b4", X"3d8af975", X"3d8b944c", X"3d8c3c76", X"3d8b48a8", X"3d8a80cc", X"3d8b459b", 
X"3d8a7103", X"3d8b87ad", X"3d8b1ee2", X"3d8a25c4", X"3d8b0555", X"3d898d9d", X"3d8acbf9", X"3d8b38ed", 
X"3d8a2b8b", X"3d89c50d", X"3d89cc82", X"3d89b3a3", X"3d8abc84", X"3d8a2791", X"3d892a26", X"3d8a37d8", 
X"3d88bf7c", X"3d89e88c", X"3d8a3108", X"3d896914", X"3d896e79", X"3d88dcc5", X"3d892a7f", X"3d89ea90", 
X"3d893a44", X"3d88afa3", X"3d89cb65", X"3d88b6b5", X"3d89adfd", X"3d89a394", X"3d88e738", X"3d89c29f", 
X"3d889e93", X"3d897557", X"3d89ef81", X"3d8919a3", X"3d88aac5", X"3d89683d", X"3d88c820", X"3d89b1f9", 
X"3d895170", X"3d88712e", X"3d897bd8", X"3d8820e9", X"3d892b6d", X"3d8993c3", X"3d889e0f", X"3d88469a", 
X"3d883cf2", X"3d886bee", X"3d895ac7", X"3d88be4c", X"3d87cf16", X"3d88dabc", X"3d8760e3", X"3d88c67a", 
X"3d88ed30", X"3d87e637", X"3d880a69", X"3d873443", X"3d87d531", X"3d889440", X"3d87c595", X"3d86f767", 
X"3d87e08a", X"3d86d065", X"3d880096", X"3d87c158", X"3d86cdc1", X"3d8798f4", X"3d863367", X"3d87109b", 
X"3d8784db", X"3d86a268", X"3d8649c6", X"3d869918", X"3d863f2d", X"3d87129d", X"3d868ed7", X"3d85c446", 
X"3d86fee5", X"3d855ed3", X"3d868de4", X"3d86b7b8", X"3d85c7d0", X"3d85f908", X"3d8579eb", X"3d85de88", 
X"3d86a0f1", X"3d85e20a", X"3d84d2d1", X"3d85f2b8", X"3d84bf09", X"3d85fde8", X"3d85dbad", X"3d84d1fb", 
X"3d8548ca", X"3d843998", X"3d854e19", X"3d85ed19", X"3d84f919", X"3d843227", X"3d84dc01", X"3d848476", 
X"3d85a33d", X"3d854862", X"3d844c93", X"3d854499", X"3d83e443", X"3d8533d3", X"3d859f91", X"3d84d1f6", 
X"3d8490b9", X"3d84b36f", X"3d84aaaa", X"3d858feb", X"3d850faa", X"3d8449a0", X"3d859f4a", X"3d8458e3", 
X"3d85813b", X"3d85ac29", X"3d84ee1e", X"3d8554a7", X"3d84bd89", X"3d857eb3", X"3d862513", X"3d856f09", 
X"3d84d015", X"3d860658", X"3d851b24", X"3d863199", X"3d860a1f", X"3d85153c", X"3d85e2de", X"3d84d228", 
X"3d85e978", X"3d8672d8", X"3d859493", X"3d84d987", X"3d858417", X"3d85244a", X"3d865432", X"3d85ee37", 
X"3d84d7dd", X"3d85d552", X"3d846a57", X"3d85cf58", X"3d86361f", X"3d85473b", X"3d85058c", X"3d84c44a", 
X"3d852356", X"3d85fe35", X"3d85640c", X"3d846f4a", X"3d8594ba", X"3d841fdc", X"3d857e19", X"3d857dca", 
X"3d847bd2", X"3d84e573", X"3d83f46d", X"3d84a2ac", X"3d85402c", X"3d847875", X"3d83a640", X"3d849239", 
X"3d83b46b", X"3d84ca4b", X"3d847d6a", X"3d83884f", X"3d847eaa", X"3d830d3a", X"3d84380e", X"3d8499a2", 
X"3d83c115", X"3d836784", X"3d838f4b", X"3d8379be", X"3d8465aa", X"3d83e0a3", X"3d82b458", X"3d83e309", 
X"3d824b4e", X"3d83ab21", X"3d83cdf9", X"3d82cffa", X"3d82ce76", X"3d82312e", X"3d82c9c2", X"3d839ff7", 
X"3d82e83a", X"3d81a904", X"3d82c3ea", X"3d81d470", X"3d832ec9", X"3d831ac2", X"3d822751", X"3d829ace", 
X"3d817a7b", X"3d829ebf", X"3d833e7e", X"3d829175", X"3d81dead", X"3d828aae", X"3d81f2f1", X"3d83005f", 
X"3d82be4e", X"3d81d24b", X"3d82ed7d", X"3d8178f6", X"3d82a68a", X"3d82ffeb", X"3d824d66", X"3d821631", 
X"3d82281b", X"3d8232c4", X"3d83106f", X"3d8295e1", X"3d81b400", X"3d82fe3d", X"3d81be8b", X"3d82f93b", 
X"3d831aa2", X"3d8240ca", X"3d826609", X"3d81b64e", X"3d82822c", X"3d833abc", X"3d82991b", X"3d818116", 
X"3d828894", X"3d816baf", X"3d82df93", X"3d82c401", X"3d81ae68", X"3d823906", X"3d80fdac", X"3d821e96", 
X"3d82bc5e", X"3d81f111", X"3d8111ed", X"3d817fb8", X"3d811f5c", X"3d823a21", X"3d81dd52", X"3d80d2f8", 
X"3d81d8de", X"3d8052f6", X"3d81a2cf", X"3d81e417", X"3d8100d8", X"3d80c9d0", X"3d806be8", X"3d809d3d", 
X"3d81674e", X"3d80dc65", X"3d7fa14e", X"3d80f320", X"3d7edf37", X"3d80b4fe", X"3d80ac7d", X"3d7f73cd", 
X"3d801e0c", X"3d7e2361", X"3d7fa056", X"3d806ba4", X"3d7f82ed", X"3d7dc390", X"3d7f66ba", X"3d7de3ad", 
X"3d80135c", X"3d7f8c7d", X"3d7d6839", X"3d7eefe8", X"3d7c0a02", X"3d7e8ae4", X"3d7f47ad", X"3d7d8512", 
X"3d7c4df1", X"3d7c73d0", X"3d7c765c", X"3d7e8f1c", X"3d7d9d14", X"3d7b1d3f", X"3d7d4e4d", X"3d7a6194", 
X"3d7d47a5", X"3d7da082", X"3d7bff8a", X"3d7bba71", X"3d7ab137", X"3d7bb454", X"3d7d6a4e", X"3d7c70e4", 
X"3d7a92a0", X"3d7c8ecf", X"3d7a6749", X"3d7cb488", X"3d7ca991", X"3d7b1cfc", X"3d7c290e", X"3d79db30", 
X"3d7bad62", X"3d7cbb9b", X"3d7b9813", X"3d7a5d53", X"3d7bd172", X"3d7a7364", X"3d7c8c0a", X"3d7c000a", 
X"3d7a2450", X"3d7c2b13", X"3d797208", X"3d7bb2b7", X"3d7c5ad9", X"3d7afdf5", X"3d7a14ba", X"3d7a3035", 
X"3d7a594b", X"3d7c410e", X"3d7b63a0", X"3d79302e", X"3d7b2549", X"3d783c16", X"3d7b0a6f", X"3d7b60b0", 
X"3d799686", X"3d797194", X"3d77f105", X"3d792c34", X"3d7ac34f", X"3d798fc7", X"3d775df5", X"3d79043f", 
X"3d76ae71", X"3d795718", X"3d79125d", X"3d773588", X"3d783e42", X"3d75b723", X"3d778a3f", X"3d789124", 
X"3d773348", X"3d75c65b", X"3d766b99", X"3d755ebf", X"3d773cbf", X"3d767f77", X"3d749ae6", X"3d766de1", 
X"3d731142", X"3d754c7b", X"3d75b0d6", X"3d74223a", X"3d73c7ec", X"3d72ee5d", X"3d731614", X"3d749cb7", 
X"3d73a1ea", X"3d719c0c", X"3d73b51d", X"3d70e9b7", X"3d7360b9", X"3d733db9", X"3d717224", X"3d71dd22", 
X"3d6fe428", X"3d715610", X"3d728732", X"3d7129f2", X"3d6f2046", X"3d705e32", X"3d6f0767", X"3d714986", 
X"3d70b1cc", X"3d6ea404", X"3d6ff02b", X"3d6d2167", X"3d6f9dd9", X"3d706958", X"3d6efdf0", X"3d6dd209", 
X"3d6e1bad", X"3d6dae84", X"3d6fa729", X"3d6efe03", X"3d6d383d", X"3d6f25f6", X"3d6c81ea", X"3d6ebdd6", 
X"3d6f1f37", X"3d6df307", X"3d6df490", X"3d6d1289", X"3d6db87d", X"3d6f1c7f", X"3d6e2e34", X"3d6cce63", 
X"3d6ecf6c", X"3d6c96cb", X"3d6ea5ff", X"3d6e837f", X"3d6d0b8f", X"3d6e1e1c", X"3d6c04c6", X"3d6dab88", 
X"3d6eaaf0", X"3d6d80af", X"3d6bffaf", X"3d6d4fcf", X"3d6c0137", X"3d6e4970", X"3d6dc63f", X"3d6be92e", 
X"3d6d597e", X"3d6adf47", X"3d6d2165", X"3d6df0f6", X"3d6c82bb", X"3d6b7719", X"3d6b58ea", X"3d6b6bfc", 
X"3d6d42e8", X"3d6c5482", X"3d6a507b", X"3d6c0fb8", X"3d692be4", X"3d6bbfce", X"3d6be7c8", X"3d6a559a", 
X"3d6a719f", X"3d690880", X"3d6a004c", X"3d6b58b5", X"3d6a3485", X"3d686b33", X"3d6a1300", X"3d67e9d8", 
X"3d6a1935", X"3d69ba63", X"3d682745", X"3d6954d5", X"3d66c1a7", X"3d685129", X"3d691c04", X"3d67d1bd", 
X"3d669dd2", X"3d671a10", X"3d66365b", X"3d67f5d6", X"3d673adb", X"3d658787", X"3d675a87", X"3d6450eb", 
X"3d66a795", X"3d66f1bc", X"3d654eee", X"3d64d662", X"3d6411c3", X"3d64879d", X"3d661c1a", X"3d65077c", 
X"3d62e27f", X"3d64d1c2", X"3d6299d3", X"3d650637", X"3d64db42", X"3d633a22", X"3d638227", X"3d61a18f", 
X"3d63485d", X"3d64879c", X"3d634d7e", X"3d61b568", X"3d62eae1", X"3d6190c8", X"3d63aaaf", X"3d635cba", 
X"3d61df84", X"3d6322b7", X"3d608d87", X"3d629068", X"3d63542b", X"3d624b7e", X"3d619a33", X"3d620a1c", 
X"3d617f5d", X"3d633a14", X"3d629051", X"3d6146fd", X"3d634ff9", X"3d60cf62", X"3d62bb37", X"3d630301", 
X"3d61e6fe", X"3d61e833", X"3d60f291", X"3d61b95f", X"3d6303a6", X"3d620d92", X"3d608828", X"3d6262db", 
X"3d60206d", X"3d628599", X"3d6266db", X"3d60d932", X"3d6166c6", X"3d5f9453", X"3d612f20", X"3d626443", 
X"3d6130bb", X"3d5fb162", X"3d60b8a7", X"3d5f8d9c", X"3d61ce3e", X"3d613cea", X"3d5f8b7a", X"3d60ca41", 
X"3d5e20b2", X"3d6032dd", X"3d60daa5", X"3d5f8bd4", X"3d5edde0", X"3d5e9638", X"3d5e94cd", X"3d602334", 
X"3d5f2ee5", X"3d5d8738", X"3d5f5b12", X"3d5c8547", X"3d5eaf2e", X"3d5eb74a", X"3d5d65a6", X"3d5dd589", 
X"3d5c445c", X"3d5d02ea", X"3d5e30e8", X"3d5d113d", X"3d5b9994", X"3d5d16a9", X"3d5b2f75", X"3d5d0876", 
X"3d5c9b68", X"3d5b444d", X"3d5c6ffe", X"3d59edae", X"3d5ba0ed", X"3d5c5d2e", X"3d5af2e4", X"3d59df01", 
X"3d5a362e", X"3d59a844", X"3d5b6b9c", X"3d5a8dca", X"3d58be11", X"3d5a83d0", X"3d57f411", X"3d5a4044", 
X"3d5a8d0d", X"3d59162b", X"3d58b95a", X"3d57f983", X"3d58aa43", X"3d5a42c2", X"3d5930d1", X"3d577cd8", 
X"3d592b7b", X"3d573beb", X"3d593832", X"3d594a0d", X"3d581b72", X"3d5896fb", X"3d56cb0c", X"3d5820a2", 
X"3d5938d0", X"3d582fd4", X"3d5733bc", X"3d588a17", X"3d571162", X"3d58d21c", X"3d587172", X"3d574923", 
X"3d58fd92", X"3d56a8bf", X"3d585cb2", X"3d59018e", X"3d57f2b2", X"3d575066", X"3d5790ae", X"3d574461", 
X"3d58c5eb", X"3d57fa19", X"3d568ef2", X"3d585834", X"3d55f158", X"3d57ffef", X"3d585818", X"3d56f11b", 
X"3d56c0f9", X"3d55cadf", X"3d569f44", X"3d580eed", X"3d56f693", X"3d556136", X"3d56f71c", X"3d54da5a", 
X"3d573c59", X"3d570842", X"3d5584ab", X"3d5631b8", X"3d543969", X"3d55a348", X"3d56a920", X"3d557274", 
X"3d543b15", X"3d54ff7f", X"3d53f77c", X"3d55b366", X"3d54fc02", X"3d537f8a", X"3d54f352", X"3d523fcb", 
X"3d540225", X"3d54798f", X"3d532cba", X"3d52d1db", X"3d524447", X"3d522456", X"3d537c41", X"3d52838d", 
X"3d51169a", X"3d52e431", X"3d505c44", X"3d523dfc", X"3d5230d5", X"3d50edeb", X"3d516dc5", X"3d4fc84b", 
X"3d50b209", X"3d51c802", X"3d508944", X"3d4efb2c", X"3d50304a", X"3d4ec3d9", X"3d508703", X"3d4ff987", 
X"3d4e7a92", X"3d4f8f75", X"3d4d4246", X"3d4f18d8", X"3d4fd15d", X"3d4e6021", X"3d4d8026", X"3d4dba31", 
X"3d4d90dc", X"3d4f4d47", X"3d4e7de0", X"3d4ced92", X"3d4ea633", X"3d4c6ea0", X"3d4e45be", X"3d4eb84f", 
X"3d4daac3", X"3d4d6eb7", X"3d4cbf3e", X"3d4d1a88", X"3d4e6e2b", X"3d4d7e52", X"3d4c6f8f", X"3d4e3125", 
X"3d4c4c72", X"3d4de451", X"3d4de0a5", X"3d4cda0b", X"3d4dd7d8", X"3d4c174f", X"3d4d5a2d", X"3d4e442d", 
X"3d4d32f3", X"3d4c6127", X"3d4d9bb6", X"3d4c76ec", X"3d4e1762", X"3d4d9899", X"3d4c54d4", X"3d4dcb81", 
X"3d4bbd30", X"3d4d50fd", X"3d4e07df", X"3d4cbd81", X"3d4bfb1d", X"3d4c1e84", X"3d4c1cd0", X"3d4daeb5", 
X"3d4ccc23", X"3d4b4b29", X"3d4ceabd", X"3d4a92f2", X"3d4cb508", X"3d4cf822", X"3d4b8bdb", X"3d4ba581", 
X"3d4a82ae", X"3d4b50d9", X"3d4c892c", X"3d4b6ef9", X"3d4a1c8a", X"3d4ba2e8", X"3d49d962", X"3d4bb385", 
X"3d4b549a", X"3d49ea82", X"3d4aeb57", X"3d48e7a8", X"3d4a220f", X"3d4aea93", X"3d49b495", X"3d48d1fe", 
X"3d4961c2", X"3d4890f2", X"3d49f75a", X"3d4936dd", X"3d47e02e", X"3d498208", X"3d4707fd", X"3d48cb0d", 
X"3d491b54", X"3d47d58a", X"3d47d710", X"3d47499a", X"3d479c12", X"3d48e174", X"3d47ce56", X"3d4620c4", 
X"3d47e142", X"3d45e3c1", X"3d47b2b2", X"3d478741", X"3d461214", X"3d468faf", X"3d451066", X"3d465773", 
X"3d4762d8", X"3d460dd1", X"3d44a38e", X"3d45b719", X"3d44eda5", X"3d46b07f", X"3d4632c4", X"3d44c48a", 
X"3d46062c", X"3d43fa91", X"3d45cdde", X"3d468d9c", X"3d4583b0", X"3d44db27", X"3d45455d", X"3d44e254", 
X"3d4651c4", X"3d45a408", X"3d447028", X"3d4651e1", X"3d444982", X"3d45d404", X"3d462305", X"3d45257b", 
X"3d4567a4", X"3d44af89", X"3d455986", X"3d467195", X"3d457be3", X"3d44694c", X"3d462349", X"3d448b4d", 
X"3d462b16", X"3d46097c", X"3d44c723", X"3d45b13e", X"3d4423c9", X"3d457a3b", X"3d467172", X"3d454642", 
X"3d440167", X"3d450c90", X"3d440edc", X"3d45e748", X"3d45623e", X"3d43e094", X"3d452841", X"3d430ff6", 
X"3d44cd25", X"3d457938", X"3d441a46", X"3d436bd9", X"3d4339ae", X"3d435cc0", X"3d44b596", X"3d43d377", 
X"3d426f10", X"3d442395", X"3d41ea35", X"3d43df88", X"3d43f00e", X"3d428928", X"3d42e7a5", X"3d41b22a", 
X"3d425ec0", X"3d435eff", X"3d425525", X"3d41024a", X"3d425bd9", X"3d40b036", X"3d423f37", X"3d41d76c", 
X"3d408902", X"3d41a160", X"3d3f8a58", X"3d40e092", X"3d4181ba", X"3d405046", X"3d3f8f68", X"3d3ff7fb", 
X"3d3f97a0", X"3d40f935", X"3d4032e0", X"3d3e9a66", X"3d404007", X"3d3e067f", X"3d3fe9be", X"3d4023c0", 
X"3d3eb336", X"3d3e822f", X"3d3de48f", X"3d3e8237", X"3d3fc4bd", X"3d3eb4aa", X"3d3cec6a", X"3d3e929a", 
X"3d3d0fb6", X"3d3eebe4", X"3d3ed3f4", X"3d3d8594", X"3d3dff3f", X"3d3c8f3e", X"3d3de47e", X"3d3ee55b", 
X"3d3ded53", X"3d3cefbc", X"3d3e1cc7", X"3d3d277c", X"3d3eab21", X"3d3e5667", X"3d3d1e8f", X"3d3ea3f7", 
X"3d3caf50", X"3d3e33a5", X"3d3ec91b", X"3d3dd154", X"3d3d6957", X"3d3dc882", X"3d3d9207", X"3d3ee4ce", 
X"3d3e2a91", X"3d3ced88", X"3d3ec1c8", X"3d3cde93", X"3d3e6b14", X"3d3ea351", X"3d3d8004", X"3d3d8fa3", 
X"3d3cdd0c", X"3d3dbdee", X"3d3edd5a", X"3d3de90f", X"3d3c7cb9", X"3d3e17c2", X"3d3c676b", X"3d3e79dc", 
X"3d3e579b", X"3d3ceb56", X"3d3d9c89", X"3d3c0c3c", X"3d3d6e0d", X"3d3e6388", X"3d3d3234", X"3d3bee8e", 
X"3d3cbb50", X"3d3bfd64", X"3d3d9b85", X"3d3d0aa0", X"3d3b97e4", X"3d3cf931", X"3d3ad117", X"3d3c8937", 
X"3d3cfa31", X"3d3bb5fe", X"3d3b51f3", X"3d3b15d0", X"3d3b3779", X"3d3c62b6", X"3d3b8e73", X"3d3a293e", 
X"3d3bcc30", X"3d398c4f", X"3d3b43b1", X"3d3b363f", X"3d39ecde", X"3d3a5bba", X"3d3904a5", X"3d39d3ec", 
X"3d3ab8f8", X"3d39bc7f", X"3d38719c", X"3d39ab59", X"3d386624", X"3d39f679", X"3d398520", X"3d380f9e", 
X"3d391604", X"3d3721fe", X"3d38c506", X"3d395b26", X"3d3815cf", X"3d3734b7", X"3d378dc1", X"3d377264", 
X"3d38dee4", X"3d381740", X"3d365f88", X"3d37f8c4", X"3d36001d", X"3d37f15a", X"3d383278", X"3d36fe0f", 
X"3d36b63f", X"3d36393d", X"3d36c32b", X"3d38023c", X"3d373515", X"3d35ecb4", X"3d377236", X"3d35e469", 
X"3d37771b", X"3d3777c1", X"3d366ae2", X"3d372902", X"3d35bf97", X"3d36f742", X"3d37ca01", X"3d36edc2", 
X"3d36253c", X"3d3758b1", X"3d364b37", X"3d37b91c", X"3d374d47", X"3d3612fa", X"3d378eae", X"3d35b0b7", 
X"3d3726da", X"3d37a787", X"3d369f4b", X"3d35ed10", X"3d36381b", X"3d3631d8", X"3d378e19", X"3d36d88d", 
X"3d356124", X"3d36ec76", X"3d34fa16", X"3d36f0e8", X"3d3732b1", X"3d35ed37", X"3d35e3fb", X"3d351122", 
X"3d35f736", X"3d3719d1", X"3d361f4b", X"3d34a294", X"3d35f4d9", X"3d344069", X"3d361669", X"3d35d976", 
X"3d34795c", X"3d353dfe", X"3d338d1a", X"3d34cd81", X"3d358af7", X"3d346d3d", X"3d3356fa", X"3d3405b5", 
X"3d335160", X"3d34a5c5", X"3d340e9a", X"3d32c36b", X"3d3423dd", X"3d31e3a8", X"3d337caa", X"3d33c66c", 
X"3d329516", X"3d3248ea", X"3d31dbcd", X"3d320114", X"3d330fb2", X"3d32416c", X"3d30dc21", X"3d3279d5", 
X"3d307de6", X"3d32342f", X"3d32158c", X"3d30bad9", X"3d310578", X"3d2fb98b", X"3d30c607", X"3d31a41d", 
X"3d308b7e", X"3d2f18ed", X"3d304123", X"3d2f5c39", X"3d30f78c", X"3d3082d3", X"3d2f0ff8", X"3d300946", 
X"3d2e31a3", X"3d2ff7cc", X"3d308c8d", X"3d2f68e4", X"3d2e8bb7", X"3d2ef0db", X"3d2ea9fb", X"3d300aef", 
X"3d2f8591", X"3d2e31a4", X"3d2fa4a5", X"3d2dc13e", X"3d2f5316", X"3d2fa271", X"3d2eb28c", X"3d2e9fe1", 
X"3d2e23c3", X"3d2e9773", X"3d2fa04c", X"3d2ee78f", X"3d2df56b", X"3d2f9711", X"3d2e0fa6", X"3d2f894a", 
X"3d2f77ef", X"3d2e67fa", X"3d2f1eb9", X"3d2db10b", X"3d2edb00", X"3d2f9052", X"3d2ea503", X"3d2d8d47", 
X"3d2eabb5", X"3d2da48f", X"3d2f407a", X"3d2ed558", X"3d2d7174", X"3d2e7f0b", X"3d2cb63e", X"3d2e4e62", 
X"3d2ee80b", X"3d2dc825", X"3d2d09ae", X"3d2d1ef9", X"3d2d31cd", X"3d2e8900", X"3d2dcf57", X"3d2c5373", 
X"3d2db2c3", X"3d2ba1bb", X"3d2d76f4", X"3d2d974c", X"3d2c5d0d", X"3d2c6858", X"3d2b70b9", X"3d2c1ea7", 
X"3d2d0c7e", X"3d2c1b63", X"3d2ab93b", X"3d2c0c52", X"3d2a6b97", X"3d2bf87f", X"3d2baa6b", X"3d2a72dd", 
X"3d2b4445", X"3d297657", X"3d2aa207", X"3d2b387f", X"3d2a30ff", X"3d294da2", X"3d29d6fa", X"3d29414f", 
X"3d2a797d", X"3d29e5f3", X"3d28a5e1", X"3d2a0847", X"3d27e595", X"3d299470", X"3d29cb5c", X"3d2888f6", 
X"3d282bea", X"3d27bcc4", X"3d280f21", X"3d292afe", X"3d28498b", X"3d26a6f6", X"3d283007", X"3d269181", 
X"3d284c39", X"3d28287e", X"3d26f10d", X"3d2737cc", X"3d260477", X"3d274c0d", X"3d2830e0", X"3d273a6c", 
X"3d2606ec", X"3d271bef", X"3d263341", X"3d27aecd", X"3d277039", X"3d264b93", X"3d274446", X"3d257b3a", 
X"3d26fa01", X"3d27895d", X"3d26aee0", X"3d261b86", X"3d269c5c", X"3d2635c6", X"3d276eb4", X"3d26eb11", 
X"3d25e366", X"3d278380", X"3d25bff8", X"3d273587", X"3d276c8e", X"3d268d49", X"3d268db1", X"3d2603c9", 
X"3d26a833", X"3d2799d0", X"3d26d802", X"3d25acd9", X"3d271fb3", X"3d258036", X"3d273d68", X"3d27277f", 
X"3d25efdc", X"3d265cac", X"3d251305", X"3d2647cd", X"3d272193", X"3d2629d9", X"3d24f55c", X"3d25c7f6", 
X"3d24d20a", X"3d26591f", X"3d25de15", X"3d247d24", X"3d253f0d", X"3d23449d", X"3d248a64", X"3d24e5b2", 
X"3d23ce7b", X"3d22f2cc", X"3d229c8c", X"3d224a1c", X"3d232ee8", X"3d2267c2", X"3d20e4c5", X"3d21c57f", 
X"3d1f7a0a", X"3d2097a1", X"3d208199", X"3d1f42ed", X"3d1ef087", X"3d1d79a8", X"3d1d6e38", X"3d1df49c", 
X"3d1d0970", X"3d1b6505", X"3d1be439", X"3d1a0a13", X"3d1aceee", X"3d1a616c", X"3d1909c2", X"3d191464", 
X"3d16e394", X"3d17451a", X"3d1784ef", X"3d164704", X"3d14a189", X"3d143acc", X"3d13013f", X"3d13a672", 
X"3d12df53", X"3d10e84c", X"3d1122de", X"3d0eaab1", X"3d0f4f01", X"3d0f3488", X"3d0db296", X"3d0c581b", 
X"3d0b1322", X"3d0a637d", X"3d0ae91f", X"3d09f354", X"3d07cae2", X"3d07f4d7", X"3d05a090", X"3d060114", 
X"3d05caaf", X"3d045c3b", X"3d0364f0", X"3d014c3f", X"3d00d4fe", X"3d01208f", X"3d0014ef", X"3cfc4dec", 
X"3cfc33f3", X"3cf7b029", X"3cf86ff7", X"3cf785cf", X"3cf468ed", X"3cf409d8", X"3cef35de", X"3cef3be2", 
X"3cef61b3", X"3ced2f62", X"3ce9fc9b", X"3ce8a299", X"3ce5e9fe", X"3ce6b4d5", X"3ce53b06", X"3ce1dd62", 
X"3ce1f04b", X"3cdd5761", X"3cddf7f7", X"3cddb76b", X"3cdb380c", X"3cd8f765", X"3cd633a8", X"3cd52cd0", 
X"3cd5ddf2", X"3cd404d2", X"3cd098a6", X"3cd0a271", X"3ccc7663", X"3ccdad97", X"3cccd64f", X"3cca2886", 
X"3cc8ff25", X"3cc53cfa", X"3cc4f27d", X"3cc53f39", X"3cc357fe", X"3cc0737e", X"3cbf96cd", X"3cbcb320", 
X"3cbd7cf8", X"3cbc2b0e", X"3cb99043", X"3cb94796", X"3cb50a4c", X"3cb568c8", X"3cb53456", X"3cb35bbb", 
X"3cb17d4e", X"3caf43e7", X"3cad98d6", X"3cae1c10", X"3cacae28", X"3caa3af8", X"3caa45eb", X"3ca66a07", 
X"3ca71859", X"3ca68084", X"3ca4ceb0", X"3ca3d62e", X"3ca0e25a", X"3ca042f8", X"3ca094a0", X"3c9f0afd", 
X"3c9c6c2c", X"3c9bf1b6", X"3c993aeb", X"3c99f63d", X"3c98f66c", X"3c970f3e", X"3c968b53", X"3c933d88", 
X"3c938a84", X"3c93847a", X"3c91edfc", X"3c90181a", X"3c8ee77a", X"3c8d7abb", X"3c8e36b5", X"3c8d11bf", 
X"3c8b28d9", X"3c8b1974", X"3c8843bb", X"3c88d4fd", X"3c889b5d", X"3c878b15", X"3c866824", X"3c84c456", 
X"3c83d397", X"3c845868", X"3c8358ef", X"3c81d765", X"3c81eae3", X"3c7ee76c", X"3c7fee00", X"3c7ed328", 
X"3c7cf1df", X"3c7c8637", X"3c77e215", X"3c77f30c", X"3c784831", X"3c7669d9", X"3c7460f6", X"3c73b75c", 
X"3c6fff0e", X"3c714e3f", X"3c6fb8e6", X"3c6d9484", X"3c6d7ee1", X"3c68a16d", X"3c692793", X"3c68cb72", 
X"3c66dd52", X"3c654011", X"3c63248e", X"3c6116e9", X"3c62279c", X"3c602622", X"3c5dc558", X"3c5e0f2f", 
X"3c593b4e", X"3c5a89d5", X"3c596a23", X"3c57402a", X"3c5684c1", X"3c52edf9", X"3c520c8d", X"3c527148", 
X"3c5021bf", X"3c4e1b65", X"3c4dc72e", X"3c49a13e", X"3c4a9aac", X"3c48b34e", X"3c4688be", X"3c4669b7", 
X"3c422291", X"3c41e713", X"3c4185b9", X"3c3f7fea", X"3c3df538", X"3c3c4211", X"3c397fc8", X"3c3a38dc", 
X"3c3813ac", X"3c3679ff", X"3c369593", X"3c31f909", X"3c3270e4", X"3c319adc", X"3c2fd591", X"3c2f29cd", 
X"3c2c6dc5", X"3c2b0011", X"3c2b64b5", X"3c292ffe", X"3c272a87", X"3c2715ee", X"3c2378a6", X"3c243ed1", 
X"3c22aaae", X"3c20ac2d", X"3c2055d1", X"3c1d2845", X"3c1c946a", X"3c1c8b57", X"3c1a39de", X"3c18739e", 
X"3c17fb06", X"3c159be0", X"3c165957", X"3c148274", X"3c12b6db", X"3c132df8", X"3c101cc6", X"3c101523", 
X"3c0fbef2", X"3c0dda75", X"3c0cf8f2", X"3c0c3780", X"3c0a3cc9", X"3c0adc11", X"3c093c80", X"3c078d54", 
X"3c080b01", X"3c051eb2", X"3c0546ad", X"3c049a37", X"3c030f07", X"3c02ce19", X"3c00fb81", X"3bff98e3", 
X"3c003589", X"3bfcd5d8", X"3bfa754a", X"3bfb4dc9", X"3bf625a8", X"3bf71719", X"3bf4dde4", X"3bf1ea0c", 
X"3bf1e9be", X"3bedb1bb", X"3bece4cd", X"3bed85aa", X"3bea4362", X"3be8443c", X"3be7c756", X"3be39d37", 
X"3be4d4bc", X"3be1c730", X"3bdf12e7", X"3bdfb583", X"3bdb077f", X"3bdad4e8", X"3bd99623", X"3bd67465", 
X"3bd50378", X"3bd2f567", X"3bcf6f93", X"3bd00c7a", X"3bcca94b", X"3bc9d86b", X"3bca6ff0", X"3bc53afe", 
X"3bc58569", X"3bc3957a", X"3bc08619", X"3bbf80a5", X"3bbc696d", X"3bbabf6e", X"3bba84b4", X"3bb7d592", 
X"3bb56a9b", X"3bb564f6", X"3bb20572", X"3bb24a70", X"3bb08076", X"3bada215", X"3bad4c7f", X"3ba9f9fd", 
X"3ba8f9da", X"3ba897fb", X"3ba5c2d7", X"3ba3a95d", X"3ba2455b", X"3b9fa296", X"3b9f76d8", X"3b9d40ac", 
X"3b9ae343", X"3b9b401d", X"3b977d24", X"3b973711", X"3b95ffea", X"3b935b14", X"3b9234a9", X"3b91649e", 
X"3b8f5f47", X"3b8fc9e5", X"3b8daca6", X"3b8af46c", X"3b8bbee1", X"3b89d415", X"3b89c144", X"3b88473b", 
X"3b866f9f", X"3b8646a4", X"3b84a257", X"3b824934", X"3b824bb1", X"3b80273b", X"3b7dd954", X"3b7f0835", 
X"3b7bec1d", X"3b7cf84d", X"3b789319", X"3b74974f", X"3b75444d", X"3b715eec", X"3b6fa21d", X"3b6ea489"
);


begin

rom_select: process (clk, en, reset)
begin
	if (rising_edge(clk)) then
			data_out <= ENVELOPE_ROM(conv_integer(index));
	end if;
end process rom_select;

end rtl;
